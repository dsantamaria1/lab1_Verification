
module fifo_DW01_mux_any_256_4_16_1 ( A, SEL, MUX );
input  [255:0] A;
input  [3:0] SEL;
output [15:0] MUX;
    wire \tmp[3][136] , \tmp[3][14] , \tmp[3][132] , \tmp[3][10] , 
        \tmp[3][139] , \tmp[3][130] , \tmp[3][129] , \tmp[3][12] , 
        \tmp[3][134] , \tmp[3][1] , \tmp[3][8] , \tmp[3][141] , \tmp[3][5] , 
        \tmp[3][7] , \tmp[3][143] , \tmp[3][3] , \tmp[3][142] , \tmp[3][2] , 
        \tmp[3][6] , \tmp[3][4] , \tmp[3][0] , \tmp[3][9] , \tmp[3][140] , 
        \tmp[3][135] , \tmp[3][138] , \tmp[3][13] , \tmp[3][131] , 
        \tmp[3][128] , \tmp[3][11] , \tmp[3][133] , \tmp[3][137] , 
        \tmp[3][15] , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
        n50, n51, n52, n56, n58, n59;
    MUX81P MX8_1_1_0 ( .D0(A[0]), .D1(A[16]), .D2(A[32]), .D3(A[48]), .D4(A
        [64]), .D5(A[80]), .D6(A[96]), .D7(A[112]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][0] ) );
    MUX81P MX8_1_1_1 ( .D0(A[1]), .D1(A[17]), .D2(A[33]), .D3(A[49]), .D4(A
        [65]), .D5(A[81]), .D6(A[97]), .D7(A[113]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][1] ) );
    MUX81P MX8_1_1_2 ( .D0(A[2]), .D1(A[18]), .D2(A[34]), .D3(A[50]), .D4(A
        [66]), .D5(A[82]), .D6(A[98]), .D7(A[114]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][2] ) );
    MUX81P MX8_1_5_10 ( .D0(A[138]), .D1(A[154]), .D2(A[170]), .D3(A[186]), 
        .D4(A[202]), .D5(A[218]), .D6(A[234]), .D7(A[250]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][138] ) );
    MUX81P MX8_1_1_3 ( .D0(A[3]), .D1(A[19]), .D2(A[35]), .D3(A[51]), .D4(A
        [67]), .D5(A[83]), .D6(A[99]), .D7(A[115]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][3] ) );
    MUX81P MX8_1_1_4 ( .D0(A[4]), .D1(A[20]), .D2(A[36]), .D3(A[52]), .D4(A
        [68]), .D5(A[84]), .D6(A[100]), .D7(A[116]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][4] ) );
    MUX81P MX8_1_1_5 ( .D0(A[5]), .D1(A[21]), .D2(A[37]), .D3(A[53]), .D4(A
        [69]), .D5(A[85]), .D6(A[101]), .D7(A[117]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][5] ) );
    MUX81P MX8_1_1_11 ( .D0(A[11]), .D1(A[27]), .D2(A[43]), .D3(A[59]), .D4(A
        [75]), .D5(A[91]), .D6(A[107]), .D7(A[123]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][11] ) );
    MUX81P MX8_1_5_3 ( .D0(A[131]), .D1(A[147]), .D2(A[163]), .D3(A[179]), 
        .D4(A[195]), .D5(A[211]), .D6(A[227]), .D7(A[243]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][131] ) );
    MUX81P MX8_1_5_4 ( .D0(A[132]), .D1(A[148]), .D2(A[164]), .D3(A[180]), 
        .D4(A[196]), .D5(A[212]), .D6(A[228]), .D7(A[244]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][132] ) );
    MUX81P MX8_1_1_10 ( .D0(A[10]), .D1(A[26]), .D2(A[42]), .D3(A[58]), .D4(A
        [74]), .D5(A[90]), .D6(A[106]), .D7(A[122]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][10] ) );
    MUX81P MX8_1_5_2 ( .D0(A[130]), .D1(A[146]), .D2(A[162]), .D3(A[178]), 
        .D4(A[194]), .D5(A[210]), .D6(A[226]), .D7(A[242]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][130] ) );
    MUX81P MX8_1_5_5 ( .D0(A[133]), .D1(A[149]), .D2(A[165]), .D3(A[181]), 
        .D4(A[197]), .D5(A[213]), .D6(A[229]), .D7(A[245]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][133] ) );
    MUX81P MX8_1_5_11 ( .D0(A[139]), .D1(A[155]), .D2(A[171]), .D3(A[187]), 
        .D4(A[203]), .D5(A[219]), .D6(A[235]), .D7(A[251]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][139] ) );
    MUX81P MX8_1_1_8 ( .D0(A[8]), .D1(A[24]), .D2(A[40]), .D3(A[56]), .D4(A
        [72]), .D5(A[88]), .D6(A[104]), .D7(A[120]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][8] ) );
    MUX81P MX8_1_5_13 ( .D0(A[141]), .D1(A[157]), .D2(A[173]), .D3(A[189]), 
        .D4(A[205]), .D5(A[221]), .D6(A[237]), .D7(A[253]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][141] ) );
    MUX81P MX8_1_1_6 ( .D0(A[6]), .D1(A[22]), .D2(A[38]), .D3(A[54]), .D4(A
        [70]), .D5(A[86]), .D6(A[102]), .D7(A[118]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][6] ) );
    MUX81P MX8_1_1_12 ( .D0(A[12]), .D1(A[28]), .D2(A[44]), .D3(A[60]), .D4(A
        [76]), .D5(A[92]), .D6(A[108]), .D7(A[124]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][12] ) );
    MUX81P MX8_1_1_15 ( .D0(A[15]), .D1(A[31]), .D2(A[47]), .D3(A[63]), .D4(A
        [79]), .D5(A[95]), .D6(A[111]), .D7(A[127]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][15] ) );
    MUX81P MX8_1_5_0 ( .D0(A[128]), .D1(A[144]), .D2(A[160]), .D3(A[176]), 
        .D4(A[192]), .D5(A[208]), .D6(A[224]), .D7(A[240]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][128] ) );
    MUX81P MX8_1_5_7 ( .D0(A[135]), .D1(A[151]), .D2(A[167]), .D3(A[183]), 
        .D4(A[199]), .D5(A[215]), .D6(A[231]), .D7(A[247]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][135] ) );
    MUX81P MX8_1_1_7 ( .D0(A[7]), .D1(A[23]), .D2(A[39]), .D3(A[55]), .D4(A
        [71]), .D5(A[87]), .D6(A[103]), .D7(A[119]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][7] ) );
    MUX81P MX8_1_5_9 ( .D0(A[137]), .D1(A[153]), .D2(A[169]), .D3(A[185]), 
        .D4(A[201]), .D5(A[217]), .D6(A[233]), .D7(A[249]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][137] ) );
    MUX81P MX8_1_5_14 ( .D0(A[142]), .D1(A[158]), .D2(A[174]), .D3(A[190]), 
        .D4(A[206]), .D5(A[222]), .D6(A[238]), .D7(A[254]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][142] ) );
    MUX81P MX8_1_1_9 ( .D0(A[9]), .D1(A[25]), .D2(A[41]), .D3(A[57]), .D4(A
        [73]), .D5(A[89]), .D6(A[105]), .D7(A[121]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][9] ) );
    MUX81P MX8_1_1_14 ( .D0(A[14]), .D1(A[30]), .D2(A[46]), .D3(A[62]), .D4(A
        [78]), .D5(A[94]), .D6(A[110]), .D7(A[126]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][14] ) );
    MUX81P MX8_1_5_1 ( .D0(A[129]), .D1(A[145]), .D2(A[161]), .D3(A[177]), 
        .D4(A[193]), .D5(A[209]), .D6(A[225]), .D7(A[241]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][129] ) );
    MUX81P MX8_1_5_8 ( .D0(A[136]), .D1(A[152]), .D2(A[168]), .D3(A[184]), 
        .D4(A[200]), .D5(A[216]), .D6(A[232]), .D7(A[248]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][136] ) );
    MUX81P MX8_1_5_15 ( .D0(A[143]), .D1(A[159]), .D2(A[175]), .D3(A[191]), 
        .D4(A[207]), .D5(A[223]), .D6(A[239]), .D7(A[255]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][143] ) );
    MUX81P MX8_1_5_12 ( .D0(A[140]), .D1(A[156]), .D2(A[172]), .D3(A[188]), 
        .D4(A[204]), .D5(A[220]), .D6(A[236]), .D7(A[252]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][140] ) );
    MUX81P MX8_1_1_13 ( .D0(A[13]), .D1(A[29]), .D2(A[45]), .D3(A[61]), .D4(A
        [77]), .D5(A[93]), .D6(A[109]), .D7(A[125]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][13] ) );
    MUX81P MX8_1_5_6 ( .D0(A[134]), .D1(A[150]), .D2(A[166]), .D3(A[182]), 
        .D4(A[198]), .D5(A[214]), .D6(A[230]), .D7(A[246]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][134] ) );
    AO2 U72 ( .A(\tmp[3][9] ), .B(n40), .C(\tmp[3][137] ), .D(SEL[3]), .Z(n39)
         );
    AO2 U73 ( .A(\tmp[3][8] ), .B(n40), .C(\tmp[3][136] ), .D(SEL[3]), .Z(n41)
         );
    AO2 U74 ( .A(\tmp[3][7] ), .B(n40), .C(\tmp[3][135] ), .D(SEL[3]), .Z(n42)
         );
    AO2 U75 ( .A(\tmp[3][6] ), .B(n40), .C(\tmp[3][134] ), .D(SEL[3]), .Z(n43)
         );
    AO2 U76 ( .A(\tmp[3][5] ), .B(n40), .C(\tmp[3][133] ), .D(SEL[3]), .Z(n44)
         );
    AO2 U77 ( .A(\tmp[3][4] ), .B(n40), .C(\tmp[3][132] ), .D(SEL[3]), .Z(n45)
         );
    AO2 U78 ( .A(\tmp[3][3] ), .B(n40), .C(\tmp[3][131] ), .D(SEL[3]), .Z(n46)
         );
    AO2 U79 ( .A(\tmp[3][2] ), .B(n40), .C(\tmp[3][130] ), .D(SEL[3]), .Z(n47)
         );
    AO2 U80 ( .A(\tmp[3][1] ), .B(n40), .C(\tmp[3][129] ), .D(SEL[3]), .Z(n48)
         );
    AO2 U81 ( .A(\tmp[3][15] ), .B(n40), .C(\tmp[3][143] ), .D(SEL[3]), .Z(n49
        ) );
    AO2 U82 ( .A(\tmp[3][14] ), .B(n40), .C(\tmp[3][142] ), .D(SEL[3]), .Z(n50
        ) );
    AO2 U83 ( .A(\tmp[3][13] ), .B(n40), .C(\tmp[3][141] ), .D(SEL[3]), .Z(n51
        ) );
    AO2 U84 ( .A(\tmp[3][12] ), .B(n40), .C(\tmp[3][140] ), .D(SEL[3]), .Z(n52
        ) );
    AO2 U85 ( .A(\tmp[3][11] ), .B(n40), .C(\tmp[3][139] ), .D(SEL[3]), .Z(n56
        ) );
    AO2 U86 ( .A(\tmp[3][10] ), .B(n40), .C(\tmp[3][138] ), .D(SEL[3]), .Z(n58
        ) );
    AO2 U87 ( .A(\tmp[3][0] ), .B(n40), .C(\tmp[3][128] ), .D(SEL[3]), .Z(n59)
         );
    IV U88 ( .A(SEL[3]), .Z(n40) );
    IV U89 ( .A(n39), .Z(MUX[9]) );
    IV U90 ( .A(n41), .Z(MUX[8]) );
    IV U91 ( .A(n42), .Z(MUX[7]) );
    IV U92 ( .A(n43), .Z(MUX[6]) );
    IV U93 ( .A(n44), .Z(MUX[5]) );
    IV U94 ( .A(n45), .Z(MUX[4]) );
    IV U95 ( .A(n46), .Z(MUX[3]) );
    IV U96 ( .A(n47), .Z(MUX[2]) );
    IV U97 ( .A(n48), .Z(MUX[1]) );
    IV U98 ( .A(n49), .Z(MUX[15]) );
    IV U99 ( .A(n50), .Z(MUX[14]) );
    IV U100 ( .A(n51), .Z(MUX[13]) );
    IV U101 ( .A(n52), .Z(MUX[12]) );
    IV U102 ( .A(n56), .Z(MUX[11]) );
    IV U103 ( .A(n58), .Z(MUX[10]) );
    IV U104 ( .A(n59), .Z(MUX[0]) );
endmodule


module fifo_DW_MEM_R_W_S_LAT_16_16_1 ( clk, wr_n, rd_addr, wr_addr, data_in, 
    data_out );
output [15:0] data_out;
input  [3:0] rd_addr;
input  [15:0] wr_addr;
input  [15:0] data_in;
input  clk, wr_n;
    wire \q[15][15] , \q[15][14] , \q[15][12] , \q[15][9] , \q[15][6] , 
        \q[15][2] , \q[14][1] , \q[10][15] , \q[6][0] , \q[1][12] , 
        \din[15][0] , \q[11][13] , \q[11][9] , \q[10][3] , \din[11][2] , 
        \din[5][1] , \din[1][3] , \q[2][2] , \din[6][12] , \q[9][14] , 
        \q[8][4] , \din[0][9] , \din[10][8] , \q[6][10] , \q[3][8] , \q[3][1] , 
        \din[10][10] , \din[8][10] , \q[0][14] , \q[11][0] , \din[10][1] , 
        \din[14][3] , \din[0][0] , \din[4][2] , \q[14][8] , \q[7][3] , 
        \din[7][14] , \din[1][10] , \q[14][5] , \q[10][7] , \q[9][10] , 
        \q[9][7] , \q[8][12] , \q[6][9] , \din[15][9] , \din[5][8] , \q[8][0] , 
        \din[10][14] , \din[8][14] , \q[2][6] , \din[11][6] , \din[0][12] , 
        \din[15][4] , \din[1][7] , \din[5][5] , \q[10][11] , \q[7][12] , 
        \q[9][3] , \q[6][4] , \din[9][12] , \q[7][7] , \din[11][12] , 
        \din[14][7] , \din[7][10] , \din[1][14] , \q[15][4] , \q[11][4] , 
        \q[8][9] , \din[10][5] , \din[4][6] , \din[0][4] , \q[7][5] , 
        \q[6][14] , \q[3][5] , \q[0][10] , \din[14][5] , \din[7][12] , 
        \din[4][4] , \q[15][0] , \q[14][7] , \q[11][15] , \q[11][6] , 
        \din[10][7] , \q[3][7] , \din[0][6] , \q[0][12] , \q[10][5] , 
        \q[9][8] , \q[9][1] , \q[8][14] , \din[11][10] , \din[9][10] , 
        \q[2][4] , \din[6][14] , \din[0][10] , \din[11][4] , \din[1][5] , 
        \din[15][6] , \q[11][11] , \q[10][13] , \q[6][6] , \din[5][7] , 
        \q[10][8] , \q[9][12] , \q[8][2] , \q[7][10] , \q[1][14] , \q[8][10] , 
        \q[2][9] , \din[11][14] , \din[9][14] , \q[9][5] , \din[1][8] , 
        \q[3][3] , \din[11][9] , \q[11][2] , \q[6][12] , \din[10][3] , 
        \din[0][2] , \din[14][1] , \q[8][6] , \q[7][1] , \din[4][0] , 
        \din[1][12] , \q[7][8] , \din[10][12] , \q[14][3] , \q[7][14] , 
        \q[1][10] , \din[14][8] , \din[8][12] , \din[4][9] , \q[6][2] , 
        \din[15][2] , \din[5][3] , \q[12][7] , \q[10][1] , \din[11][0] , 
        \q[4][4] , \q[2][0] , \din[1][1] , \wren[8] , \din[6][10] , 
        \din[0][14] , \din[5][11] , \din[3][15] , \din[7][5] , \q[0][6] , 
        \din[13][6] , \din[3][7] , \q[14][14] , \q[13][4] , \q[4][15] , 
        \q[2][11] , \q[1][5] , \din[13][13] , \din[9][1] , \din[2][13] , 
        \din[9][8] , \din[2][4] , \q[12][10] , \q[5][13] , \din[12][5] , 
        \din[6][6] , \q[14][12] , \q[14][10] , \q[13][12] , \q[13][9] , 
        \q[5][7] , \q[1][8] , \wren[1] , \din[14][11] , \din[12][15] , 
        \din[15][13] , \din[8][2] , \din[12][8] , \din[9][5] , \q[4][11] , 
        \q[2][15] , \din[2][9] , \q[12][3] , \q[0][2] , \din[3][3] , \q[4][9] , 
        \q[4][0] , \din[13][2] , \din[7][1] , \din[8][6] , \din[5][15] , 
        \din[3][11] , \wren[5] , \din[14][15] , \din[12][11] , \din[7][8] , 
        \q[13][0] , \q[12][14] , \q[5][3] , \q[3][13] , \din[6][2] , 
        \q[5][15] , \q[1][1] , \wren[13] , \din[2][0] , \din[12][1] , 
        \din[4][13] , \q[3][11] , \q[13][10] , \q[13][2] , \q[5][1] , 
        \wren[11] , \din[6][0] , \din[2][2] , \q[12][8] , \q[1][3] , 
        \din[12][3] , \din[4][11] , \din[2][15] , \din[13][9] , \q[0][9] , 
        \din[3][8] , \q[0][0] , \wren[7] , \din[12][13] , \din[8][4] , 
        \q[15][11] , \q[15][10] , \q[13][6] , \q[12][1] , \q[4][13] , 
        \q[5][8] , \q[4][2] , \din[13][0] , \din[3][1] , \din[7][3] , 
        \din[3][13] , \din[6][9] , \q[1][7] , \wren[3] , \din[15][11] , 
        \din[9][7] , \din[13][15] , \din[14][13] , \din[8][0] , \din[4][15] , 
        \din[2][11] , \q[12][12] , \wren[15] , \din[2][6] , \din[12][7] , 
        \din[6][4] , \q[12][5] , \q[5][11] , \q[3][15] , \q[5][5] , \q[4][6] , 
        \din[15][15] , \din[13][11] , \din[9][3] , \din[7][7] , \din[5][13] , 
        \din[3][5] , \q[2][13] , \din[13][4] , \q[13][15] , \q[13][14] , 
        \q[13][7] , \q[0][4] , \wren[14] , \wren[2] , \din[8][9] , 
        \din[14][12] , \din[8][1] , \q[12][13] , \q[1][6] , \din[12][6] , 
        \din[2][7] , \din[4][14] , \din[2][10] , \q[5][10] , \q[5][4] , 
        \q[3][14] , \q[4][7] , \din[15][14] , \din[6][5] , \din[13][10] , 
        \din[9][2] , \din[7][6] , \din[5][12] , \q[2][12] , \q[0][5] , 
        \din[8][8] , \q[14][13] , \q[12][4] , \din[3][4] , \q[5][14] , 
        \q[3][10] , \din[13][5] , \din[6][1] , \q[13][3] , \q[5][0] , 
        \q[1][2] , \din[4][10] , \din[2][14] , \din[2][3] , \q[12][9] , 
        \q[0][8] , \wren[10] , \din[12][2] , \din[8][5] , \din[13][8] , 
        \q[12][0] , \wren[6] , \din[12][12] , \din[3][9] , \din[13][1] , 
        \din[3][0] , \q[15][13] , \q[14][11] , \q[13][13] , \q[13][11] , 
        \q[13][8] , \q[5][9] , \q[4][12] , \q[4][3] , \q[0][1] , \din[7][2] , 
        \din[3][12] , \din[15][10] , \din[13][14] , \din[9][6] , \din[6][8] , 
        \din[12][9] , \q[12][2] , \q[1][9] , \din[15][12] , \din[2][8] , 
        \din[9][4] , \din[3][2] , \q[4][10] , \q[0][3] , \din[13][3] , 
        \q[2][14] , \q[12][15] , \q[4][8] , \q[4][1] , \din[5][14] , 
        \din[3][10] , \din[8][7] , \din[7][0] , \din[7][9] , \wren[4] , 
        \din[14][14] , \din[12][10] , \din[6][3] , \q[13][1] , \q[5][2] , 
        \q[3][12] , \q[1][0] , \din[4][12] , \wren[12] , \q[4][5] , \wren[9] , 
        \din[12][0] , \din[2][1] , \din[7][4] , \din[5][10] , \din[3][14] , 
        \q[15][8] , \q[15][1] , \q[14][15] , \q[13][5] , \q[12][6] , 
        \q[4][14] , \q[2][10] , \q[0][7] , \din[13][12] , \din[13][7] , 
        \din[3][6] , \din[9][0] , \din[2][5] , \q[5][12] , \q[1][4] , 
        \din[12][4] , \din[9][9] , \din[2][12] , \q[12][11] , \q[11][10] , 
        \q[11][3] , \q[10][9] , \q[8][11] , \q[5][6] , \din[6][7] , \wren[0] , 
        \din[14][10] , \din[12][14] , \din[8][3] , \q[9][4] , \din[9][15] , 
        \q[2][8] , \din[11][15] , \din[11][8] , \din[1][9] , \din[10][2] , 
        \din[0][3] , \q[3][2] , \q[7][0] , \q[6][13] , \din[14][0] , 
        \din[1][13] , \q[8][7] , \din[4][1] , \q[15][7] , \q[15][5] , 
        \q[14][2] , \q[7][9] , \din[14][9] , \din[8][13] , \din[4][8] , 
        \din[10][13] , \din[15][3] , \din[5][2] , \q[10][0] , \q[7][15] , 
        \q[6][3] , \q[2][1] , \q[1][11] , \din[6][11] , \din[0][15] , 
        \din[11][1] , \din[14][4] , \din[1][0] , \din[4][5] , \q[14][6] , 
        \q[11][14] , \q[7][4] , \q[3][6] , \din[7][13] , \q[0][13] , 
        \q[11][7] , \din[10][6] , \q[10][12] , \q[10][4] , \q[9][9] , 
        \q[9][0] , \din[11][11] , \din[0][7] , \q[8][15] , \din[9][11] , 
        \din[11][5] , \din[1][4] , \q[2][5] , \din[6][15] , \din[0][11] , 
        \q[7][11] , \q[1][15] , \q[6][7] , \din[15][7] , \q[14][4] , 
        \q[10][10] , \q[10][6] , \q[9][13] , \q[8][3] , \din[5][6] , 
        \q[9][11] , \q[8][1] , \din[10][15] , \din[8][15] , \din[11][7] , 
        \q[7][13] , \q[6][5] , \q[2][7] , \din[1][6] , \din[0][13] , 
        \din[15][5] , \din[5][4] , \q[9][2] , \din[11][13] , \din[9][13] , 
        \din[14][6] , \q[15][3] , \q[14][0] , \q[11][5] , \q[8][8] , \q[7][6] , 
        \din[4][7] , \q[6][15] , \q[3][4] , \din[7][11] , \din[1][15] , 
        \q[0][11] , \din[10][4] , \din[0][5] , \din[15][1] , \q[11][12] , 
        \q[11][8] , \q[10][14] , \din[5][0] , \q[10][2] , \q[6][1] , 
        \q[1][13] , \q[2][3] , \din[11][3] , \din[6][13] , \din[1][2] , 
        \q[3][9] , \q[11][1] , \q[9][15] , \q[8][5] , \din[0][8] , 
        \din[10][11] , \din[10][9] , \din[8][11] , \din[10][0] , \q[6][11] , 
        \q[3][0] , \din[0][1] , \q[0][15] , \q[7][2] , \din[14][2] , 
        \din[7][15] , \din[1][11] , \din[4][3] , \q[14][9] , \q[6][8] , 
        \q[9][6] , \q[8][13] , \din[15][8] , \din[5][9] , n38, n60, n61, n62, 
        n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n108, n109;
    fifo_DW01_mux_any_256_4_16_1 MX ( .A({\q[15][15] , \q[15][14] , 
        \q[15][13] , \q[15][12] , \q[15][11] , \q[15][10] , \q[15][9] , 
        \q[15][8] , \q[15][7] , \q[15][6] , \q[15][5] , \q[15][4] , \q[15][3] , 
        \q[15][2] , \q[15][1] , \q[15][0] , \q[14][15] , \q[14][14] , 
        \q[14][13] , \q[14][12] , \q[14][11] , \q[14][10] , \q[14][9] , 
        \q[14][8] , \q[14][7] , \q[14][6] , \q[14][5] , \q[14][4] , \q[14][3] , 
        \q[14][2] , \q[14][1] , \q[14][0] , \q[13][15] , \q[13][14] , 
        \q[13][13] , \q[13][12] , \q[13][11] , \q[13][10] , \q[13][9] , 
        \q[13][8] , \q[13][7] , \q[13][6] , \q[13][5] , \q[13][4] , \q[13][3] , 
        \q[13][2] , \q[13][1] , \q[13][0] , \q[12][15] , \q[12][14] , 
        \q[12][13] , \q[12][12] , \q[12][11] , \q[12][10] , \q[12][9] , 
        \q[12][8] , \q[12][7] , \q[12][6] , \q[12][5] , \q[12][4] , \q[12][3] , 
        \q[12][2] , \q[12][1] , \q[12][0] , \q[11][15] , \q[11][14] , 
        \q[11][13] , \q[11][12] , \q[11][11] , \q[11][10] , \q[11][9] , 
        \q[11][8] , \q[11][7] , \q[11][6] , \q[11][5] , \q[11][4] , \q[11][3] , 
        \q[11][2] , \q[11][1] , \q[11][0] , \q[10][15] , \q[10][14] , 
        \q[10][13] , \q[10][12] , \q[10][11] , \q[10][10] , \q[10][9] , 
        \q[10][8] , \q[10][7] , \q[10][6] , \q[10][5] , \q[10][4] , \q[10][3] , 
        \q[10][2] , \q[10][1] , \q[10][0] , \q[9][15] , \q[9][14] , \q[9][13] , 
        \q[9][12] , \q[9][11] , \q[9][10] , \q[9][9] , \q[9][8] , \q[9][7] , 
        \q[9][6] , \q[9][5] , \q[9][4] , \q[9][3] , \q[9][2] , \q[9][1] , 
        \q[9][0] , \q[8][15] , \q[8][14] , \q[8][13] , \q[8][12] , \q[8][11] , 
        \q[8][10] , \q[8][9] , \q[8][8] , \q[8][7] , \q[8][6] , \q[8][5] , 
        \q[8][4] , \q[8][3] , \q[8][2] , \q[8][1] , \q[8][0] , \q[7][15] , 
        \q[7][14] , \q[7][13] , \q[7][12] , \q[7][11] , \q[7][10] , \q[7][9] , 
        \q[7][8] , \q[7][7] , \q[7][6] , \q[7][5] , \q[7][4] , \q[7][3] , 
        \q[7][2] , \q[7][1] , \q[7][0] , \q[6][15] , \q[6][14] , \q[6][13] , 
        \q[6][12] , \q[6][11] , \q[6][10] , \q[6][9] , \q[6][8] , \q[6][7] , 
        \q[6][6] , \q[6][5] , \q[6][4] , \q[6][3] , \q[6][2] , \q[6][1] , 
        \q[6][0] , \q[5][15] , \q[5][14] , \q[5][13] , \q[5][12] , \q[5][11] , 
        \q[5][10] , \q[5][9] , \q[5][8] , \q[5][7] , \q[5][6] , \q[5][5] , 
        \q[5][4] , \q[5][3] , \q[5][2] , \q[5][1] , \q[5][0] , \q[4][15] , 
        \q[4][14] , \q[4][13] , \q[4][12] , \q[4][11] , \q[4][10] , \q[4][9] , 
        \q[4][8] , \q[4][7] , \q[4][6] , \q[4][5] , \q[4][4] , \q[4][3] , 
        \q[4][2] , \q[4][1] , \q[4][0] , \q[3][15] , \q[3][14] , \q[3][13] , 
        \q[3][12] , \q[3][11] , \q[3][10] , \q[3][9] , \q[3][8] , \q[3][7] , 
        \q[3][6] , \q[3][5] , \q[3][4] , \q[3][3] , \q[3][2] , \q[3][1] , 
        \q[3][0] , \q[2][15] , \q[2][14] , \q[2][13] , \q[2][12] , \q[2][11] , 
        \q[2][10] , \q[2][9] , \q[2][8] , \q[2][7] , \q[2][6] , \q[2][5] , 
        \q[2][4] , \q[2][3] , \q[2][2] , \q[2][1] , \q[2][0] , \q[1][15] , 
        \q[1][14] , \q[1][13] , \q[1][12] , \q[1][11] , \q[1][10] , \q[1][9] , 
        \q[1][8] , \q[1][7] , \q[1][6] , \q[1][5] , \q[1][4] , \q[1][3] , 
        \q[1][2] , \q[1][1] , \q[1][0] , \q[0][15] , \q[0][14] , \q[0][13] , 
        \q[0][12] , \q[0][11] , \q[0][10] , \q[0][9] , \q[0][8] , \q[0][7] , 
        \q[0][6] , \q[0][5] , \q[0][4] , \q[0][3] , \q[0][2] , \q[0][1] , 
        \q[0][0] }), .SEL(rd_addr), .MUX(data_out) );
    MUX21H MX1_0_0 ( .A(\q[0][0] ), .B(data_in[0]), .S(\wren[0] ), .Z(
        \din[0][0] ) );
    MUX21H MX1_0_11 ( .A(\q[11][0] ), .B(data_in[0]), .S(\wren[11] ), .Z(
        \din[11][0] ) );
    MUX21H MX1_8_1 ( .A(\q[1][8] ), .B(data_in[8]), .S(\wren[1] ), .Z(
        \din[1][8] ) );
    MUX21H MX1_15_9 ( .A(\q[9][15] ), .B(data_in[15]), .S(\wren[9] ), .Z(
        \din[9][15] ) );
    MUX21H MX1_12_3 ( .A(\q[3][12] ), .B(data_in[12]), .S(\wren[3] ), .Z(
        \din[3][12] ) );
    MUX21H MX1_14_12 ( .A(\q[12][14] ), .B(data_in[14]), .S(\wren[12] ), .Z(
        \din[12][14] ) );
    MUX21H MX1_5_6 ( .A(\q[6][5] ), .B(data_in[5]), .S(\wren[6] ), .Z(
        \din[6][5] ) );
    MUX21H MX1_6_14 ( .A(\q[14][6] ), .B(data_in[6]), .S(\wren[14] ), .Z(
        \din[14][6] ) );
    MUX21H MX1_1_0 ( .A(\q[0][1] ), .B(data_in[1]), .S(\wren[0] ), .Z(
        \din[0][1] ) );
    MUX21H MX1_4_6 ( .A(\q[6][4] ), .B(data_in[4]), .S(\wren[6] ), .Z(
        \din[6][4] ) );
    MUX21H MX1_1_10 ( .A(\q[10][1] ), .B(data_in[1]), .S(\wren[10] ), .Z(
        \din[10][1] ) );
    MUX21H MX1_0_9 ( .A(\q[9][0] ), .B(data_in[0]), .S(\wren[9] ), .Z(
        \din[9][0] ) );
    MUX21H MX1_4_10 ( .A(\q[10][4] ), .B(data_in[4]), .S(\wren[10] ), .Z(
        \din[10][4] ) );
    MUX21H MX1_14_9 ( .A(\q[9][14] ), .B(data_in[14]), .S(\wren[9] ), .Z(
        \din[9][14] ) );
    MUX21H MX1_7_15 ( .A(\q[15][7] ), .B(data_in[7]), .S(\wren[15] ), .Z(
        \din[15][7] ) );
    MUX21H MX1_15_13 ( .A(\q[13][15] ), .B(data_in[15]), .S(\wren[13] ), .Z(
        \din[13][15] ) );
    MUX21H MX1_9_1 ( .A(\q[1][9] ), .B(data_in[9]), .S(\wren[1] ), .Z(
        \din[1][9] ) );
    MUX21H MX1_8_8 ( .A(\q[8][8] ), .B(data_in[8]), .S(\wren[8] ), .Z(
        \din[8][8] ) );
    MUX21H MX1_13_3 ( .A(\q[3][13] ), .B(data_in[13]), .S(\wren[3] ), .Z(
        \din[3][13] ) );
    MUX21H MX1_15_0 ( .A(\q[0][15] ), .B(data_in[15]), .S(\wren[0] ), .Z(
        \din[0][15] ) );
    MUX21H MX1_10_6 ( .A(\q[6][10] ), .B(data_in[10]), .S(\wren[6] ), .Z(
        \din[6][10] ) );
    MUX21H MX1_1_9 ( .A(\q[9][1] ), .B(data_in[1]), .S(\wren[9] ), .Z(
        \din[9][1] ) );
    MUX21H MX1_2_5 ( .A(\q[5][2] ), .B(data_in[2]), .S(\wren[5] ), .Z(
        \din[5][2] ) );
    MUX21H MX1_8_13 ( .A(\q[13][8] ), .B(data_in[8]), .S(\wren[13] ), .Z(
        \din[13][8] ) );
    MUX21H MX1_2_15 ( .A(\q[15][2] ), .B(data_in[2]), .S(\wren[15] ), .Z(
        \din[15][2] ) );
    MUX21H MX1_7_3 ( .A(\q[3][7] ), .B(data_in[7]), .S(\wren[3] ), .Z(
        \din[3][7] ) );
    MUX21H MX1_10_13 ( .A(\q[13][10] ), .B(data_in[10]), .S(\wren[13] ), .Z(
        \din[13][10] ) );
    MUX21H MX1_5_11 ( .A(\q[11][5] ), .B(data_in[5]), .S(\wren[11] ), .Z(
        \din[11][5] ) );
    MUX21H MX1_6_3 ( .A(\q[3][6] ), .B(data_in[6]), .S(\wren[3] ), .Z(
        \din[3][6] ) );
    MUX21H MX1_3_5 ( .A(\q[5][3] ), .B(data_in[3]), .S(\wren[5] ), .Z(
        \din[5][3] ) );
    MUX21H MX1_3_14 ( .A(\q[14][3] ), .B(data_in[3]), .S(\wren[14] ), .Z(
        \din[14][3] ) );
    MUX21H MX1_9_8 ( .A(\q[8][9] ), .B(data_in[9]), .S(\wren[8] ), .Z(
        \din[8][9] ) );
    MUX21H MX1_9_12 ( .A(\q[12][9] ), .B(data_in[9]), .S(\wren[12] ), .Z(
        \din[12][9] ) );
    MUX21H MX1_11_6 ( .A(\q[6][11] ), .B(data_in[11]), .S(\wren[6] ), .Z(
        \din[6][11] ) );
    MUX21H MX1_14_0 ( .A(\q[0][14] ), .B(data_in[14]), .S(\wren[0] ), .Z(
        \din[0][14] ) );
    MUX21H MX1_9_15 ( .A(\q[15][9] ), .B(data_in[9]), .S(\wren[15] ), .Z(
        \din[15][9] ) );
    MUX21H MX1_11_12 ( .A(\q[12][11] ), .B(data_in[11]), .S(\wren[12] ), .Z(
        \din[12][11] ) );
    MUX21H MX1_14_7 ( .A(\q[7][14] ), .B(data_in[14]), .S(\wren[7] ), .Z(
        \din[7][14] ) );
    MUX21H MX1_11_1 ( .A(\q[1][11] ), .B(data_in[11]), .S(\wren[1] ), .Z(
        \din[1][11] ) );
    MUX21H MX1_3_13 ( .A(\q[13][3] ), .B(data_in[3]), .S(\wren[13] ), .Z(
        \din[13][3] ) );
    MUX21H MX1_11_15 ( .A(\q[15][11] ), .B(data_in[11]), .S(\wren[15] ), .Z(
        \din[15][11] ) );
    MUX21H MX1_4_8 ( .A(\q[8][4] ), .B(data_in[4]), .S(\wren[8] ), .Z(
        \din[8][4] ) );
    MUX21H MX1_3_2 ( .A(\q[2][3] ), .B(data_in[3]), .S(\wren[2] ), .Z(
        \din[2][3] ) );
    MUX21H MX1_6_4 ( .A(\q[4][6] ), .B(data_in[6]), .S(\wren[4] ), .Z(
        \din[4][6] ) );
    MUX21H MX1_2_2 ( .A(\q[2][2] ), .B(data_in[2]), .S(\wren[2] ), .Z(
        \din[2][2] ) );
    MUX21H MX1_2_12 ( .A(\q[12][2] ), .B(data_in[2]), .S(\wren[12] ), .Z(
        \din[12][2] ) );
    MUX21H MX1_5_8 ( .A(\q[8][5] ), .B(data_in[5]), .S(\wren[8] ), .Z(
        \din[8][5] ) );
    MUX21H MX1_8_14 ( .A(\q[14][8] ), .B(data_in[8]), .S(\wren[14] ), .Z(
        \din[14][8] ) );
    MUX21H MX1_10_14 ( .A(\q[14][10] ), .B(data_in[10]), .S(\wren[14] ), .Z(
        \din[14][10] ) );
    MUX21H MX1_7_4 ( .A(\q[4][7] ), .B(data_in[7]), .S(\wren[4] ), .Z(
        \din[4][7] ) );
    MUX21H MX1_7_12 ( .A(\q[12][7] ), .B(data_in[7]), .S(\wren[12] ), .Z(
        \din[12][7] ) );
    MUX21H MX1_10_1 ( .A(\q[1][10] ), .B(data_in[10]), .S(\wren[1] ), .Z(
        \din[1][10] ) );
    MUX21H MX1_15_7 ( .A(\q[7][15] ), .B(data_in[15]), .S(\wren[7] ), .Z(
        \din[7][15] ) );
    MUX21H MX1_9_6 ( .A(\q[6][9] ), .B(data_in[9]), .S(\wren[6] ), .Z(
        \din[6][9] ) );
    MUX21H MX1_11_8 ( .A(\q[8][11] ), .B(data_in[11]), .S(\wren[8] ), .Z(
        \din[8][11] ) );
    MUX21H MX1_13_4 ( .A(\q[4][13] ), .B(data_in[13]), .S(\wren[4] ), .Z(
        \din[4][13] ) );
    MUX21H MX1_15_14 ( .A(\q[14][15] ), .B(data_in[15]), .S(\wren[14] ), .Z(
        \din[14][15] ) );
    MUX21H MX1_0_1 ( .A(\q[1][0] ), .B(data_in[0]), .S(\wren[1] ), .Z(
        \din[1][0] ) );
    MUX21H MX1_0_6 ( .A(\q[6][0] ), .B(data_in[0]), .S(\wren[6] ), .Z(
        \din[6][0] ) );
    MUX21H MX1_0_7 ( .A(\q[7][0] ), .B(data_in[0]), .S(\wren[7] ), .Z(
        \din[7][0] ) );
    MUX21H MX1_1_7 ( .A(\q[7][1] ), .B(data_in[1]), .S(\wren[7] ), .Z(
        \din[7][1] ) );
    MUX21H MX1_4_1 ( .A(\q[1][4] ), .B(data_in[4]), .S(\wren[1] ), .Z(
        \din[1][4] ) );
    MUX21H MX1_13_11 ( .A(\q[11][13] ), .B(data_in[13]), .S(\wren[11] ), .Z(
        \din[11][13] ) );
    MUX21H MX1_5_1 ( .A(\q[1][5] ), .B(data_in[5]), .S(\wren[1] ), .Z(
        \din[1][5] ) );
    MUX21H MX1_6_13 ( .A(\q[13][6] ), .B(data_in[6]), .S(\wren[13] ), .Z(
        \din[13][6] ) );
    MUX21H MX1_14_15 ( .A(\q[15][14] ), .B(data_in[14]), .S(\wren[15] ), .Z(
        \din[15][14] ) );
    MUX21H MX1_8_6 ( .A(\q[6][8] ), .B(data_in[8]), .S(\wren[6] ), .Z(
        \din[6][8] ) );
    MUX21H MX1_8_15 ( .A(\q[15][8] ), .B(data_in[8]), .S(\wren[15] ), .Z(
        \din[15][8] ) );
    MUX21H MX1_10_8 ( .A(\q[8][10] ), .B(data_in[10]), .S(\wren[8] ), .Z(
        \din[8][10] ) );
    MUX21H MX1_12_10 ( .A(\q[10][12] ), .B(data_in[12]), .S(\wren[10] ), .Z(
        \din[10][12] ) );
    MUX21H MX1_12_4 ( .A(\q[4][12] ), .B(data_in[12]), .S(\wren[4] ), .Z(
        \din[4][12] ) );
    MUX21H MX1_10_0 ( .A(\q[0][10] ), .B(data_in[10]), .S(\wren[0] ), .Z(
        \din[0][10] ) );
    MUX21H MX1_15_6 ( .A(\q[6][15] ), .B(data_in[15]), .S(\wren[6] ), .Z(
        \din[6][15] ) );
    MUX21H MX1_2_3 ( .A(\q[3][2] ), .B(data_in[2]), .S(\wren[3] ), .Z(
        \din[3][2] ) );
    MUX21H MX1_2_13 ( .A(\q[13][2] ), .B(data_in[2]), .S(\wren[13] ), .Z(
        \din[13][2] ) );
    MUX21H MX1_5_9 ( .A(\q[9][5] ), .B(data_in[5]), .S(\wren[9] ), .Z(
        \din[9][5] ) );
    MUX21H MX1_7_5 ( .A(\q[5][7] ), .B(data_in[7]), .S(\wren[5] ), .Z(
        \din[5][7] ) );
    MUX21H MX1_10_15 ( .A(\q[15][10] ), .B(data_in[10]), .S(\wren[15] ), .Z(
        \din[15][10] ) );
    MUX21H MX1_4_9 ( .A(\q[9][4] ), .B(data_in[4]), .S(\wren[9] ), .Z(
        \din[9][4] ) );
    MUX21H MX1_3_3 ( .A(\q[3][3] ), .B(data_in[3]), .S(\wren[3] ), .Z(
        \din[3][3] ) );
    MUX21H MX1_6_5 ( .A(\q[5][6] ), .B(data_in[6]), .S(\wren[5] ), .Z(
        \din[5][6] ) );
    MUX21H MX1_9_14 ( .A(\q[14][9] ), .B(data_in[9]), .S(\wren[14] ), .Z(
        \din[14][9] ) );
    MUX21H MX1_14_6 ( .A(\q[6][14] ), .B(data_in[14]), .S(\wren[6] ), .Z(
        \din[6][14] ) );
    MUX21H MX1_11_0 ( .A(\q[0][11] ), .B(data_in[11]), .S(\wren[0] ), .Z(
        \din[0][11] ) );
    MUX21H MX1_3_12 ( .A(\q[12][3] ), .B(data_in[3]), .S(\wren[12] ), .Z(
        \din[12][3] ) );
    MUX21H MX1_11_14 ( .A(\q[14][11] ), .B(data_in[11]), .S(\wren[14] ), .Z(
        \din[14][11] ) );
    MUX21H MX1_5_0 ( .A(\q[0][5] ), .B(data_in[5]), .S(\wren[0] ), .Z(
        \din[0][5] ) );
    MUX21H MX1_8_7 ( .A(\q[7][8] ), .B(data_in[8]), .S(\wren[7] ), .Z(
        \din[7][8] ) );
    MUX21H MX1_10_9 ( .A(\q[9][10] ), .B(data_in[10]), .S(\wren[9] ), .Z(
        \din[9][10] ) );
    MUX21H MX1_12_11 ( .A(\q[11][12] ), .B(data_in[12]), .S(\wren[11] ), .Z(
        \din[11][12] ) );
    MUX21H MX1_12_5 ( .A(\q[5][12] ), .B(data_in[12]), .S(\wren[5] ), .Z(
        \din[5][12] ) );
    MUX21H MX1_6_12 ( .A(\q[12][6] ), .B(data_in[6]), .S(\wren[12] ), .Z(
        \din[12][6] ) );
    MUX21H MX1_14_14 ( .A(\q[14][14] ), .B(data_in[14]), .S(\wren[14] ), .Z(
        \din[14][14] ) );
    MUX21H MX1_1_6 ( .A(\q[6][1] ), .B(data_in[1]), .S(\wren[6] ), .Z(
        \din[6][1] ) );
    MUX21H MX1_4_0 ( .A(\q[0][4] ), .B(data_in[4]), .S(\wren[0] ), .Z(
        \din[0][4] ) );
    MUX21H MX1_7_13 ( .A(\q[13][7] ), .B(data_in[7]), .S(\wren[13] ), .Z(
        \din[13][7] ) );
    MUX21H MX1_13_10 ( .A(\q[10][13] ), .B(data_in[13]), .S(\wren[10] ), .Z(
        \din[10][13] ) );
    MUX21H MX1_11_9 ( .A(\q[9][11] ), .B(data_in[11]), .S(\wren[9] ), .Z(
        \din[9][11] ) );
    MUX21H MX1_9_7 ( .A(\q[7][9] ), .B(data_in[9]), .S(\wren[7] ), .Z(
        \din[7][9] ) );
    MUX21H MX1_13_5 ( .A(\q[5][13] ), .B(data_in[13]), .S(\wren[5] ), .Z(
        \din[5][13] ) );
    MUX21H MX1_15_15 ( .A(\q[15][15] ), .B(data_in[15]), .S(\wren[15] ), .Z(
        \din[15][15] ) );
    MUX21H MX1_7_14 ( .A(\q[14][7] ), .B(data_in[7]), .S(\wren[14] ), .Z(
        \din[14][7] ) );
    MUX21H MX1_9_0 ( .A(\q[0][9] ), .B(data_in[9]), .S(\wren[0] ), .Z(
        \din[0][9] ) );
    MUX21H MX1_14_8 ( .A(\q[8][14] ), .B(data_in[14]), .S(\wren[8] ), .Z(
        \din[8][14] ) );
    MUX21H MX1_15_12 ( .A(\q[12][15] ), .B(data_in[15]), .S(\wren[12] ), .Z(
        \din[12][15] ) );
    MUX21H MX1_13_2 ( .A(\q[2][13] ), .B(data_in[13]), .S(\wren[2] ), .Z(
        \din[2][13] ) );
    MUX21H MX1_1_1 ( .A(\q[1][1] ), .B(data_in[1]), .S(\wren[1] ), .Z(
        \din[1][1] ) );
    MUX21H MX1_1_11 ( .A(\q[11][1] ), .B(data_in[1]), .S(\wren[11] ), .Z(
        \din[11][1] ) );
    MUX21H MX1_4_7 ( .A(\q[7][4] ), .B(data_in[4]), .S(\wren[7] ), .Z(
        \din[7][4] ) );
    MUX21H MX1_14_13 ( .A(\q[13][14] ), .B(data_in[14]), .S(\wren[13] ), .Z(
        \din[13][14] ) );
    MUX21H MX1_0_2 ( .A(\q[2][0] ), .B(data_in[0]), .S(\wren[2] ), .Z(
        \din[2][0] ) );
    MUX21H MX1_0_3 ( .A(\q[3][0] ), .B(data_in[0]), .S(\wren[3] ), .Z(
        \din[3][0] ) );
    MUX21H MX1_0_8 ( .A(\q[8][0] ), .B(data_in[0]), .S(\wren[8] ), .Z(
        \din[8][0] ) );
    MUX21H MX1_0_10 ( .A(\q[10][0] ), .B(data_in[0]), .S(\wren[10] ), .Z(
        \din[10][0] ) );
    MUX21H MX1_5_7 ( .A(\q[7][5] ), .B(data_in[5]), .S(\wren[7] ), .Z(
        \din[7][5] ) );
    MUX21H MX1_6_15 ( .A(\q[15][6] ), .B(data_in[6]), .S(\wren[15] ), .Z(
        \din[15][6] ) );
    MUX21H MX1_8_0 ( .A(\q[0][8] ), .B(data_in[8]), .S(\wren[0] ), .Z(
        \din[0][8] ) );
    MUX21H MX1_1_8 ( .A(\q[8][1] ), .B(data_in[1]), .S(\wren[8] ), .Z(
        \din[8][1] ) );
    MUX21H MX1_3_15 ( .A(\q[15][3] ), .B(data_in[3]), .S(\wren[15] ), .Z(
        \din[15][3] ) );
    MUX21H MX1_12_2 ( .A(\q[2][12] ), .B(data_in[12]), .S(\wren[2] ), .Z(
        \din[2][12] ) );
    MUX21H MX1_15_8 ( .A(\q[8][15] ), .B(data_in[15]), .S(\wren[8] ), .Z(
        \din[8][15] ) );
    MUX21H MX1_9_9 ( .A(\q[9][9] ), .B(data_in[9]), .S(\wren[9] ), .Z(
        \din[9][9] ) );
    MUX21H MX1_11_7 ( .A(\q[7][11] ), .B(data_in[11]), .S(\wren[7] ), .Z(
        \din[7][11] ) );
    MUX21H MX1_9_13 ( .A(\q[13][9] ), .B(data_in[9]), .S(\wren[13] ), .Z(
        \din[13][9] ) );
    MUX21H MX1_14_1 ( .A(\q[1][14] ), .B(data_in[14]), .S(\wren[1] ), .Z(
        \din[1][14] ) );
    MUX21H MX1_11_13 ( .A(\q[13][11] ), .B(data_in[11]), .S(\wren[13] ), .Z(
        \din[13][11] ) );
    MUX21H MX1_5_10 ( .A(\q[10][5] ), .B(data_in[5]), .S(\wren[10] ), .Z(
        \din[10][5] ) );
    MUX21H MX1_6_2 ( .A(\q[2][6] ), .B(data_in[6]), .S(\wren[2] ), .Z(
        \din[2][6] ) );
    MUX21H MX1_3_4 ( .A(\q[4][3] ), .B(data_in[3]), .S(\wren[4] ), .Z(
        \din[4][3] ) );
    MUX21H MX1_0_12 ( .A(\q[12][0] ), .B(data_in[0]), .S(\wren[12] ), .Z(
        \din[12][0] ) );
    MUX21H MX1_2_4 ( .A(\q[4][2] ), .B(data_in[2]), .S(\wren[4] ), .Z(
        \din[4][2] ) );
    MUX21H MX1_8_12 ( .A(\q[12][8] ), .B(data_in[8]), .S(\wren[12] ), .Z(
        \din[12][8] ) );
    MUX21H MX1_2_14 ( .A(\q[14][2] ), .B(data_in[2]), .S(\wren[14] ), .Z(
        \din[14][2] ) );
    MUX21H MX1_7_2 ( .A(\q[2][7] ), .B(data_in[7]), .S(\wren[2] ), .Z(
        \din[2][7] ) );
    MUX21H MX1_4_11 ( .A(\q[11][4] ), .B(data_in[4]), .S(\wren[11] ), .Z(
        \din[11][4] ) );
    MUX21H MX1_10_12 ( .A(\q[12][10] ), .B(data_in[10]), .S(\wren[12] ), .Z(
        \din[12][10] ) );
    MUX21H MX1_8_9 ( .A(\q[9][8] ), .B(data_in[8]), .S(\wren[9] ), .Z(
        \din[9][8] ) );
    MUX21H MX1_10_7 ( .A(\q[7][10] ), .B(data_in[10]), .S(\wren[7] ), .Z(
        \din[7][10] ) );
    MUX21H MX1_15_1 ( .A(\q[1][15] ), .B(data_in[15]), .S(\wren[1] ), .Z(
        \din[1][15] ) );
    MUX21H MX1_12_0 ( .A(\q[0][12] ), .B(data_in[12]), .S(\wren[0] ), .Z(
        \din[0][12] ) );
    MUX21H MX1_8_2 ( .A(\q[2][8] ), .B(data_in[8]), .S(\wren[2] ), .Z(
        \din[2][8] ) );
    MUX21H MX1_12_14 ( .A(\q[14][12] ), .B(data_in[12]), .S(\wren[14] ), .Z(
        \din[14][12] ) );
    MUX21H MX1_7_9 ( .A(\q[9][7] ), .B(data_in[7]), .S(\wren[9] ), .Z(
        \din[9][7] ) );
    MUX21H MX1_5_5 ( .A(\q[5][5] ), .B(data_in[5]), .S(\wren[5] ), .Z(
        \din[5][5] ) );
    MUX21H MX1_1_3 ( .A(\q[3][1] ), .B(data_in[1]), .S(\wren[3] ), .Z(
        \din[3][1] ) );
    MUX21H MX1_6_9 ( .A(\q[9][6] ), .B(data_in[6]), .S(\wren[9] ), .Z(
        \din[9][6] ) );
    MUX21H MX1_14_11 ( .A(\q[11][14] ), .B(data_in[14]), .S(\wren[11] ), .Z(
        \din[11][14] ) );
    MUX21H MX1_1_13 ( .A(\q[13][1] ), .B(data_in[1]), .S(\wren[13] ), .Z(
        \din[13][1] ) );
    MUX21H MX1_2_1 ( .A(\q[1][2] ), .B(data_in[2]), .S(\wren[1] ), .Z(
        \din[1][2] ) );
    MUX21H MX1_2_6 ( .A(\q[6][2] ), .B(data_in[2]), .S(\wren[6] ), .Z(
        \din[6][2] ) );
    MUX21H MX1_4_5 ( .A(\q[5][4] ), .B(data_in[4]), .S(\wren[5] ), .Z(
        \din[5][4] ) );
    MUX21H MX1_13_15 ( .A(\q[15][13] ), .B(data_in[13]), .S(\wren[15] ), .Z(
        \din[15][13] ) );
    MUX21H MX1_4_13 ( .A(\q[13][4] ), .B(data_in[4]), .S(\wren[13] ), .Z(
        \din[13][4] ) );
    MUX21H MX1_9_2 ( .A(\q[2][9] ), .B(data_in[9]), .S(\wren[2] ), .Z(
        \din[2][9] ) );
    MUX21H MX1_13_0 ( .A(\q[0][13] ), .B(data_in[13]), .S(\wren[0] ), .Z(
        \din[0][13] ) );
    MUX21H MX1_15_10 ( .A(\q[10][15] ), .B(data_in[15]), .S(\wren[10] ), .Z(
        \din[10][15] ) );
    MUX21H MX1_12_9 ( .A(\q[9][12] ), .B(data_in[12]), .S(\wren[9] ), .Z(
        \din[9][12] ) );
    MUX21H MX1_7_0 ( .A(\q[0][7] ), .B(data_in[7]), .S(\wren[0] ), .Z(
        \din[0][7] ) );
    MUX21H MX1_10_5 ( .A(\q[5][10] ), .B(data_in[10]), .S(\wren[5] ), .Z(
        \din[5][10] ) );
    MUX21H MX1_15_3 ( .A(\q[3][15] ), .B(data_in[15]), .S(\wren[3] ), .Z(
        \din[3][15] ) );
    MUX21H MX1_10_10 ( .A(\q[10][10] ), .B(data_in[10]), .S(\wren[10] ), .Z(
        \din[10][10] ) );
    MUX21H MX1_8_10 ( .A(\q[10][8] ), .B(data_in[8]), .S(\wren[10] ), .Z(
        \din[10][8] ) );
    MUX21H MX1_3_6 ( .A(\q[6][3] ), .B(data_in[3]), .S(\wren[6] ), .Z(
        \din[6][3] ) );
    MUX21H MX1_3_10 ( .A(\q[10][3] ), .B(data_in[3]), .S(\wren[10] ), .Z(
        \din[10][3] ) );
    MUX21H MX1_5_12 ( .A(\q[12][5] ), .B(data_in[5]), .S(\wren[12] ), .Z(
        \din[12][5] ) );
    MUX21H MX1_6_0 ( .A(\q[0][6] ), .B(data_in[6]), .S(\wren[0] ), .Z(
        \din[0][6] ) );
    MUX21H MX1_9_11 ( .A(\q[11][9] ), .B(data_in[9]), .S(\wren[11] ), .Z(
        \din[11][9] ) );
    MUX21H MX1_11_11 ( .A(\q[11][11] ), .B(data_in[11]), .S(\wren[11] ), .Z(
        \din[11][11] ) );
    MUX21H MX1_13_9 ( .A(\q[9][13] ), .B(data_in[13]), .S(\wren[9] ), .Z(
        \din[9][13] ) );
    MUX21H MX1_14_3 ( .A(\q[3][14] ), .B(data_in[14]), .S(\wren[3] ), .Z(
        \din[3][14] ) );
    MUX21H MX1_11_5 ( .A(\q[5][11] ), .B(data_in[11]), .S(\wren[5] ), .Z(
        \din[5][11] ) );
    MUX21H MX1_3_1 ( .A(\q[1][3] ), .B(data_in[3]), .S(\wren[1] ), .Z(
        \din[1][3] ) );
    MUX21H MX1_5_15 ( .A(\q[15][5] ), .B(data_in[5]), .S(\wren[15] ), .Z(
        \din[15][5] ) );
    MUX21H MX1_6_7 ( .A(\q[7][6] ), .B(data_in[6]), .S(\wren[7] ), .Z(
        \din[7][6] ) );
    MUX21H MX1_11_2 ( .A(\q[2][11] ), .B(data_in[11]), .S(\wren[2] ), .Z(
        \din[2][11] ) );
    MUX21H MX1_14_4 ( .A(\q[4][14] ), .B(data_in[14]), .S(\wren[4] ), .Z(
        \din[4][14] ) );
    MUX21H MX1_2_11 ( .A(\q[11][2] ), .B(data_in[2]), .S(\wren[11] ), .Z(
        \din[11][2] ) );
    MUX21H MX1_3_8 ( .A(\q[8][3] ), .B(data_in[3]), .S(\wren[8] ), .Z(
        \din[8][3] ) );
    MUX21H MX1_4_14 ( .A(\q[14][4] ), .B(data_in[4]), .S(\wren[14] ), .Z(
        \din[14][4] ) );
    MUX21H MX1_7_7 ( .A(\q[7][7] ), .B(data_in[7]), .S(\wren[7] ), .Z(
        \din[7][7] ) );
    MUX21H MX1_10_2 ( .A(\q[2][10] ), .B(data_in[10]), .S(\wren[2] ), .Z(
        \din[2][10] ) );
    MUX21H MX1_15_4 ( .A(\q[4][15] ), .B(data_in[15]), .S(\wren[4] ), .Z(
        \din[4][15] ) );
    MUX21H MX1_13_7 ( .A(\q[7][13] ), .B(data_in[13]), .S(\wren[7] ), .Z(
        \din[7][13] ) );
    MUX21H MX1_7_11 ( .A(\q[11][7] ), .B(data_in[7]), .S(\wren[11] ), .Z(
        \din[11][7] ) );
    MUX21H MX1_9_5 ( .A(\q[5][9] ), .B(data_in[9]), .S(\wren[5] ), .Z(
        \din[5][9] ) );
    MUX21H MX1_4_2 ( .A(\q[2][4] ), .B(data_in[4]), .S(\wren[2] ), .Z(
        \din[2][4] ) );
    MUX21H MX1_13_12 ( .A(\q[12][13] ), .B(data_in[13]), .S(\wren[12] ), .Z(
        \din[12][13] ) );
    MUX21H MX1_0_4 ( .A(\q[4][0] ), .B(data_in[0]), .S(\wren[4] ), .Z(
        \din[4][0] ) );
    MUX21H MX1_1_4 ( .A(\q[4][1] ), .B(data_in[1]), .S(\wren[4] ), .Z(
        \din[4][1] ) );
    MUX21H MX1_1_14 ( .A(\q[14][1] ), .B(data_in[1]), .S(\wren[14] ), .Z(
        \din[14][1] ) );
    MUX21H MX1_2_8 ( .A(\q[8][2] ), .B(data_in[2]), .S(\wren[8] ), .Z(
        \din[8][2] ) );
    MUX21H MX1_0_5 ( .A(\q[5][0] ), .B(data_in[0]), .S(\wren[5] ), .Z(
        \din[5][0] ) );
    MUX21H MX1_0_14 ( .A(\q[14][0] ), .B(data_in[0]), .S(\wren[14] ), .Z(
        \din[14][0] ) );
    MUX21H MX1_0_15 ( .A(\q[15][0] ), .B(data_in[0]), .S(\wren[15] ), .Z(
        \din[15][0] ) );
    MUX21H MX1_5_2 ( .A(\q[2][5] ), .B(data_in[5]), .S(\wren[2] ), .Z(
        \din[2][5] ) );
    MUX21H MX1_6_10 ( .A(\q[10][6] ), .B(data_in[6]), .S(\wren[10] ), .Z(
        \din[10][6] ) );
    MUX21H MX1_8_5 ( .A(\q[5][8] ), .B(data_in[8]), .S(\wren[5] ), .Z(
        \din[5][8] ) );
    MUX21H MX1_12_7 ( .A(\q[7][12] ), .B(data_in[12]), .S(\wren[7] ), .Z(
        \din[7][12] ) );
    MUX21H MX1_12_13 ( .A(\q[13][12] ), .B(data_in[12]), .S(\wren[13] ), .Z(
        \din[13][12] ) );
    MUX21H MX1_2_0 ( .A(\q[0][2] ), .B(data_in[2]), .S(\wren[0] ), .Z(
        \din[0][2] ) );
    MUX21H MX1_2_10 ( .A(\q[10][2] ), .B(data_in[2]), .S(\wren[10] ), .Z(
        \din[10][2] ) );
    MUX21H MX1_4_15 ( .A(\q[15][4] ), .B(data_in[4]), .S(\wren[15] ), .Z(
        \din[15][4] ) );
    MUX21H MX1_10_3 ( .A(\q[3][10] ), .B(data_in[10]), .S(\wren[3] ), .Z(
        \din[3][10] ) );
    MUX21H MX1_15_5 ( .A(\q[5][15] ), .B(data_in[15]), .S(\wren[5] ), .Z(
        \din[5][15] ) );
    MUX21H MX1_3_0 ( .A(\q[0][3] ), .B(data_in[3]), .S(\wren[0] ), .Z(
        \din[0][3] ) );
    MUX21H MX1_5_14 ( .A(\q[14][5] ), .B(data_in[5]), .S(\wren[14] ), .Z(
        \din[14][5] ) );
    MUX21H MX1_6_6 ( .A(\q[6][6] ), .B(data_in[6]), .S(\wren[6] ), .Z(
        \din[6][6] ) );
    MUX21H MX1_7_6 ( .A(\q[6][7] ), .B(data_in[7]), .S(\wren[6] ), .Z(
        \din[6][7] ) );
    MUX21H MX1_3_11 ( .A(\q[11][3] ), .B(data_in[3]), .S(\wren[11] ), .Z(
        \din[11][3] ) );
    MUX21H MX1_11_3 ( .A(\q[3][11] ), .B(data_in[11]), .S(\wren[3] ), .Z(
        \din[3][11] ) );
    MUX21H MX1_12_6 ( .A(\q[6][12] ), .B(data_in[12]), .S(\wren[6] ), .Z(
        \din[6][12] ) );
    MUX21H MX1_14_5 ( .A(\q[5][14] ), .B(data_in[14]), .S(\wren[5] ), .Z(
        \din[5][14] ) );
    MUX21H MX1_8_4 ( .A(\q[4][8] ), .B(data_in[8]), .S(\wren[4] ), .Z(
        \din[4][8] ) );
    MUX21H MX1_12_12 ( .A(\q[12][12] ), .B(data_in[12]), .S(\wren[12] ), .Z(
        \din[12][12] ) );
    MUX21H MX1_2_9 ( .A(\q[9][2] ), .B(data_in[2]), .S(\wren[9] ), .Z(
        \din[9][2] ) );
    MUX21H MX1_3_9 ( .A(\q[9][3] ), .B(data_in[3]), .S(\wren[9] ), .Z(
        \din[9][3] ) );
    MUX21H MX1_5_3 ( .A(\q[3][5] ), .B(data_in[5]), .S(\wren[3] ), .Z(
        \din[3][5] ) );
    MUX21H MX1_6_11 ( .A(\q[11][6] ), .B(data_in[6]), .S(\wren[11] ), .Z(
        \din[11][6] ) );
    MUX21H MX1_4_3 ( .A(\q[3][4] ), .B(data_in[4]), .S(\wren[3] ), .Z(
        \din[3][4] ) );
    MUX21H MX1_13_13 ( .A(\q[13][13] ), .B(data_in[13]), .S(\wren[13] ), .Z(
        \din[13][13] ) );
    MUX21H MX1_1_2 ( .A(\q[2][1] ), .B(data_in[1]), .S(\wren[2] ), .Z(
        \din[2][1] ) );
    MUX21H MX1_1_5 ( .A(\q[5][1] ), .B(data_in[1]), .S(\wren[5] ), .Z(
        \din[5][1] ) );
    MUX21H MX1_1_12 ( .A(\q[12][1] ), .B(data_in[1]), .S(\wren[12] ), .Z(
        \din[12][1] ) );
    MUX21H MX1_1_15 ( .A(\q[15][1] ), .B(data_in[1]), .S(\wren[15] ), .Z(
        \din[15][1] ) );
    MUX21H MX1_6_8 ( .A(\q[8][6] ), .B(data_in[6]), .S(\wren[8] ), .Z(
        \din[8][6] ) );
    MUX21H MX1_13_6 ( .A(\q[6][13] ), .B(data_in[13]), .S(\wren[6] ), .Z(
        \din[6][13] ) );
    MUX21H MX1_7_10 ( .A(\q[10][7] ), .B(data_in[7]), .S(\wren[10] ), .Z(
        \din[10][7] ) );
    MUX21H MX1_9_3 ( .A(\q[3][9] ), .B(data_in[9]), .S(\wren[3] ), .Z(
        \din[3][9] ) );
    MUX21H MX1_9_4 ( .A(\q[4][9] ), .B(data_in[9]), .S(\wren[4] ), .Z(
        \din[4][9] ) );
    MUX21H MX1_13_1 ( .A(\q[1][13] ), .B(data_in[13]), .S(\wren[1] ), .Z(
        \din[1][13] ) );
    MUX21H MX1_15_11 ( .A(\q[11][15] ), .B(data_in[15]), .S(\wren[11] ), .Z(
        \din[11][15] ) );
    MUX21H MX1_4_4 ( .A(\q[4][4] ), .B(data_in[4]), .S(\wren[4] ), .Z(
        \din[4][4] ) );
    MUX21H MX1_13_14 ( .A(\q[14][13] ), .B(data_in[13]), .S(\wren[14] ), .Z(
        \din[14][13] ) );
    MUX21H MX1_7_8 ( .A(\q[8][7] ), .B(data_in[7]), .S(\wren[8] ), .Z(
        \din[8][7] ) );
    MUX21H MX1_5_4 ( .A(\q[4][5] ), .B(data_in[5]), .S(\wren[4] ), .Z(
        \din[4][5] ) );
    MUX21H MX1_14_10 ( .A(\q[10][14] ), .B(data_in[14]), .S(\wren[10] ), .Z(
        \din[10][14] ) );
    MUX21H MX1_0_13 ( .A(\q[13][0] ), .B(data_in[0]), .S(\wren[13] ), .Z(
        \din[13][0] ) );
    MUX21H MX1_12_1 ( .A(\q[1][12] ), .B(data_in[12]), .S(\wren[1] ), .Z(
        \din[1][12] ) );
    MUX21H MX1_8_3 ( .A(\q[3][8] ), .B(data_in[8]), .S(\wren[3] ), .Z(
        \din[3][8] ) );
    MUX21H MX1_9_10 ( .A(\q[10][9] ), .B(data_in[9]), .S(\wren[10] ), .Z(
        \din[10][9] ) );
    MUX21H MX1_11_10 ( .A(\q[10][11] ), .B(data_in[11]), .S(\wren[10] ), .Z(
        \din[10][11] ) );
    MUX21H MX1_12_15 ( .A(\q[15][12] ), .B(data_in[12]), .S(\wren[15] ), .Z(
        \din[15][12] ) );
    MUX21H MX1_13_8 ( .A(\q[8][13] ), .B(data_in[13]), .S(\wren[8] ), .Z(
        \din[8][13] ) );
    MUX21H MX1_14_2 ( .A(\q[2][14] ), .B(data_in[14]), .S(\wren[2] ), .Z(
        \din[2][14] ) );
    MUX21H MX1_11_4 ( .A(\q[4][11] ), .B(data_in[11]), .S(\wren[4] ), .Z(
        \din[4][11] ) );
    MUX21H MX1_2_7 ( .A(\q[7][2] ), .B(data_in[2]), .S(\wren[7] ), .Z(
        \din[7][2] ) );
    MUX21H MX1_3_7 ( .A(\q[7][3] ), .B(data_in[3]), .S(\wren[7] ), .Z(
        \din[7][3] ) );
    MUX21H MX1_5_13 ( .A(\q[13][5] ), .B(data_in[5]), .S(\wren[13] ), .Z(
        \din[13][5] ) );
    MUX21H MX1_6_1 ( .A(\q[1][6] ), .B(data_in[6]), .S(\wren[1] ), .Z(
        \din[1][6] ) );
    MUX21H MX1_7_1 ( .A(\q[1][7] ), .B(data_in[7]), .S(\wren[1] ), .Z(
        \din[1][7] ) );
    MUX21H MX1_10_11 ( .A(\q[11][10] ), .B(data_in[10]), .S(\wren[11] ), .Z(
        \din[11][10] ) );
    MUX21H MX1_4_12 ( .A(\q[12][4] ), .B(data_in[4]), .S(\wren[12] ), .Z(
        \din[12][4] ) );
    MUX21H MX1_8_11 ( .A(\q[11][8] ), .B(data_in[8]), .S(\wren[11] ), .Z(
        \din[11][8] ) );
    MUX21H MX1_12_8 ( .A(\q[8][12] ), .B(data_in[12]), .S(\wren[8] ), .Z(
        \din[8][12] ) );
    MUX21H MX1_10_4 ( .A(\q[4][10] ), .B(data_in[10]), .S(\wren[4] ), .Z(
        \din[4][10] ) );
    MUX21H MX1_15_2 ( .A(\q[2][15] ), .B(data_in[15]), .S(\wren[2] ), .Z(
        \din[2][15] ) );
    LD1 F0_11_13 ( .D(\din[13][11] ), .G(n38), .Q(\q[13][11] ) );
    LD1 F0_14_2 ( .D(\din[2][14] ), .G(n38), .Q(\q[2][14] ) );
    LD1 F0_9_10 ( .D(\din[10][9] ), .G(n38), .Q(\q[10][9] ) );
    LD1 F0_11_4 ( .D(\din[4][11] ), .G(n38), .Q(\q[4][11] ) );
    LD1 F0_5_13 ( .D(\din[13][5] ), .G(n38), .Q(\q[13][5] ) );
    LD1 F0_3_0 ( .D(\din[0][3] ), .G(n38), .Q(\q[0][3] ) );
    LD1 F0_13_8 ( .D(\din[8][13] ), .G(n38), .Q(\q[8][13] ) );
    LD1 F0_15_2 ( .D(\din[2][15] ), .G(n38), .Q(\q[2][15] ) );
    LD1 F0_10_4 ( .D(\din[4][10] ), .G(n38), .Q(\q[4][10] ) );
    LD1 F0_6_6 ( .D(\din[6][6] ), .G(n38), .Q(\q[6][6] ) );
    LD1 F0_10_12 ( .D(\din[12][10] ), .G(n38), .Q(\q[12][10] ) );
    LD1 F0_7_6 ( .D(\din[6][7] ), .G(n38), .Q(\q[6][7] ) );
    LD1 F0_12_8 ( .D(\din[8][12] ), .G(n38), .Q(\q[8][12] ) );
    LD1 F0_8_11 ( .D(\din[11][8] ), .G(n38), .Q(\q[11][8] ) );
    LD1 F0_4_12 ( .D(\din[12][4] ), .G(n38), .Q(\q[12][4] ) );
    LD1 F0_2_0 ( .D(\din[0][2] ), .G(n38), .Q(\q[0][2] ) );
    LD1 F0_9_4 ( .D(\din[4][9] ), .G(n38), .Q(\q[4][9] ) );
    LD1 F0_1_12 ( .D(\din[12][1] ), .G(n38), .Q(\q[12][1] ) );
    LD1 F0_15_12 ( .D(\din[12][15] ), .G(n38), .Q(\q[12][15] ) );
    LD1 F0_13_1 ( .D(\din[1][13] ), .G(n38), .Q(\q[1][13] ) );
    LD1 F0_4_3 ( .D(\din[3][4] ), .G(n38), .Q(\q[3][4] ) );
    LD1 F0_5_3 ( .D(\din[3][5] ), .G(n38), .Q(\q[3][5] ) );
    LD1 F0_3_9 ( .D(\din[9][3] ), .G(n38), .Q(\q[9][3] ) );
    LD1 F0_1_5 ( .D(\din[5][1] ), .G(n38), .Q(\q[5][1] ) );
    LD1 F0_0_13 ( .D(\din[13][0] ), .G(n38), .Q(\q[13][0] ) );
    LD1 F0_14_13 ( .D(\din[13][14] ), .G(n38), .Q(\q[13][14] ) );
    LD1 F0_12_1 ( .D(\din[1][12] ), .G(n38), .Q(\q[1][12] ) );
    LD1 F0_8_4 ( .D(\din[4][8] ), .G(n38), .Q(\q[4][8] ) );
    LD1 F0_12_11 ( .D(\din[11][12] ), .G(n38), .Q(\q[11][12] ) );
    LD1 F0_8_3 ( .D(\din[3][8] ), .G(n38), .Q(\q[3][8] ) );
    LD1 F0_6_11 ( .D(\din[11][6] ), .G(n38), .Q(\q[11][6] ) );
    LD1 F0_2_9 ( .D(\din[9][2] ), .G(n38), .Q(\q[9][2] ) );
    LD1 F0_14_14 ( .D(\din[14][14] ), .G(n38), .Q(\q[14][14] ) );
    LD1 F0_0_5 ( .D(\din[5][0] ), .G(n38), .Q(\q[5][0] ) );
    LD1 F0_7_8 ( .D(\din[8][7] ), .G(n38), .Q(\q[8][7] ) );
    LD1 F0_5_4 ( .D(\din[4][5] ), .G(n38), .Q(\q[4][5] ) );
    LD1 F0_13_10 ( .D(\din[10][13] ), .G(n38), .Q(\q[10][13] ) );
    LD1 F0_12_6 ( .D(\din[6][12] ), .G(n38), .Q(\q[6][12] ) );
    LD1 F0_4_4 ( .D(\din[4][4] ), .G(n38), .Q(\q[4][4] ) );
    LD1 F0_7_10 ( .D(\din[10][7] ), .G(n38), .Q(\q[10][7] ) );
    LD1 F0_1_2 ( .D(\din[2][1] ), .G(n38), .Q(\q[2][1] ) );
    LD1 F0_0_14 ( .D(\din[14][0] ), .G(n38), .Q(\q[14][0] ) );
    LD1 F0_13_6 ( .D(\din[6][13] ), .G(n38), .Q(\q[6][13] ) );
    LD1 F0_15_15 ( .D(\din[15][15] ), .G(n38), .Q(\q[15][15] ) );
    LD1 F0_6_8 ( .D(\din[8][6] ), .G(n38), .Q(\q[8][6] ) );
    LD1 F0_9_3 ( .D(\din[3][9] ), .G(n38), .Q(\q[3][9] ) );
    LD1 F0_15_5 ( .D(\din[5][15] ), .G(n38), .Q(\q[5][15] ) );
    LD1 F0_10_3 ( .D(\din[3][10] ), .G(n38), .Q(\q[3][10] ) );
    LD1 F0_4_15 ( .D(\din[15][4] ), .G(n38), .Q(\q[15][4] ) );
    LD1 F0_2_10 ( .D(\din[10][2] ), .G(n38), .Q(\q[10][2] ) );
    LD1 F0_10_15 ( .D(\din[15][10] ), .G(n38), .Q(\q[15][10] ) );
    LD1 F0_7_1 ( .D(\din[1][7] ), .G(n38), .Q(\q[1][7] ) );
    LD1 F0_14_5 ( .D(\din[5][14] ), .G(n38), .Q(\q[5][14] ) );
    LD1 F0_11_3 ( .D(\din[3][11] ), .G(n38), .Q(\q[3][11] ) );
    LD1 F0_6_1 ( .D(\din[1][6] ), .G(n38), .Q(\q[1][6] ) );
    LD1 F0_3_11 ( .D(\din[11][3] ), .G(n38), .Q(\q[11][3] ) );
    LD1 F0_2_7 ( .D(\din[7][2] ), .G(n38), .Q(\q[7][2] ) );
    LD1 F0_11_14 ( .D(\din[14][11] ), .G(n38), .Q(\q[14][11] ) );
    LD1 F0_5_14 ( .D(\din[14][5] ), .G(n38), .Q(\q[14][5] ) );
    LD1 F0_15_14 ( .D(\din[14][15] ), .G(n38), .Q(\q[14][15] ) );
    LD1 F0_3_7 ( .D(\din[7][3] ), .G(n38), .Q(\q[7][3] ) );
    LD1 F0_1_15 ( .D(\din[15][1] ), .G(n38), .Q(\q[15][1] ) );
    LD1 F0_9_2 ( .D(\din[2][9] ), .G(n38), .Q(\q[2][9] ) );
    LD1 F0_13_11 ( .D(\din[11][13] ), .G(n38), .Q(\q[11][13] ) );
    LD1 F0_4_5 ( .D(\din[5][4] ), .G(n38), .Q(\q[5][4] ) );
    LD1 F0_1_14 ( .D(\din[14][1] ), .G(n38), .Q(\q[14][1] ) );
    LD1 F0_1_3 ( .D(\din[3][1] ), .G(n38), .Q(\q[3][1] ) );
    LD1 F0_13_7 ( .D(\din[7][13] ), .G(n38), .Q(\q[7][13] ) );
    LD1 F0_7_11 ( .D(\din[11][7] ), .G(n38), .Q(\q[11][7] ) );
    LD1 F0_6_9 ( .D(\din[9][6] ), .G(n38), .Q(\q[9][6] ) );
    LD1 F0_14_15 ( .D(\din[15][14] ), .G(n38), .Q(\q[15][14] ) );
    LD1 F0_12_7 ( .D(\din[7][12] ), .G(n38), .Q(\q[7][12] ) );
    LD1 F0_7_9 ( .D(\din[9][7] ), .G(n38), .Q(\q[9][7] ) );
    LD1 F0_5_5 ( .D(\din[5][5] ), .G(n38), .Q(\q[5][5] ) );
    LD1 F0_12_10 ( .D(\din[10][12] ), .G(n38), .Q(\q[10][12] ) );
    LD1 F0_8_2 ( .D(\din[2][8] ), .G(n38), .Q(\q[2][8] ) );
    LD1 F0_6_10 ( .D(\din[10][6] ), .G(n38), .Q(\q[10][6] ) );
    LD1 F0_11_15 ( .D(\din[15][11] ), .G(n38), .Q(\q[15][11] ) );
    LD1 F0_5_15 ( .D(\din[15][5] ), .G(n38), .Q(\q[15][5] ) );
    LD1 F0_14_4 ( .D(\din[4][14] ), .G(n38), .Q(\q[4][14] ) );
    LD1 F0_11_2 ( .D(\din[2][11] ), .G(n38), .Q(\q[2][11] ) );
    LD1 F0_6_0 ( .D(\din[0][6] ), .G(n38), .Q(\q[0][6] ) );
    LD1 F0_3_10 ( .D(\din[10][3] ), .G(n38), .Q(\q[10][3] ) );
    LD1 F0_3_6 ( .D(\din[6][3] ), .G(n38), .Q(\q[6][3] ) );
    LD1 F0_15_4 ( .D(\din[4][15] ), .G(n38), .Q(\q[4][15] ) );
    LD1 F0_10_2 ( .D(\din[2][10] ), .G(n38), .Q(\q[2][10] ) );
    LD1 F0_4_14 ( .D(\din[14][4] ), .G(n38), .Q(\q[14][4] ) );
    LD1 F0_7_0 ( .D(\din[0][7] ), .G(n38), .Q(\q[0][7] ) );
    LD1 F0_10_14 ( .D(\din[14][10] ), .G(n38), .Q(\q[14][10] ) );
    LD1 F0_15_3 ( .D(\din[3][15] ), .G(n38), .Q(\q[3][15] ) );
    LD1 F0_10_13 ( .D(\din[13][10] ), .G(n38), .Q(\q[13][10] ) );
    LD1 F0_10_5 ( .D(\din[5][10] ), .G(n38), .Q(\q[5][10] ) );
    LD1 F0_8_10 ( .D(\din[10][8] ), .G(n38), .Q(\q[10][8] ) );
    LD1 F0_12_9 ( .D(\din[9][12] ), .G(n38), .Q(\q[9][12] ) );
    LD1 F0_7_7 ( .D(\din[7][7] ), .G(n38), .Q(\q[7][7] ) );
    LD1 F0_2_11 ( .D(\din[11][2] ), .G(n38), .Q(\q[11][2] ) );
    LD1 F0_2_6 ( .D(\din[6][2] ), .G(n38), .Q(\q[6][2] ) );
    LD1 F0_14_3 ( .D(\din[3][14] ), .G(n38), .Q(\q[3][14] ) );
    LD1 F0_9_11 ( .D(\din[11][9] ), .G(n38), .Q(\q[11][9] ) );
    LD1 F0_11_5 ( .D(\din[5][11] ), .G(n38), .Q(\q[5][11] ) );
    LD1 F0_4_13 ( .D(\din[13][4] ), .G(n38), .Q(\q[13][4] ) );
    LD1 F0_13_9 ( .D(\din[9][13] ), .G(n38), .Q(\q[9][13] ) );
    LD1 F0_3_1 ( .D(\din[1][3] ), .G(n38), .Q(\q[1][3] ) );
    LD1 F0_6_7 ( .D(\din[7][6] ), .G(n38), .Q(\q[7][6] ) );
    LD1 F0_11_12 ( .D(\din[12][11] ), .G(n38), .Q(\q[12][11] ) );
    LD1 F0_8_5 ( .D(\din[5][8] ), .G(n38), .Q(\q[5][8] ) );
    LD1 F0_5_12 ( .D(\din[12][5] ), .G(n38), .Q(\q[12][5] ) );
    LD1 F0_5_2 ( .D(\din[2][5] ), .G(n38), .Q(\q[2][5] ) );
    LD1 F0_2_1 ( .D(\din[1][2] ), .G(n38), .Q(\q[1][2] ) );
    LD1 F0_0_15 ( .D(\din[15][0] ), .G(n38), .Q(\q[15][0] ) );
    LD1 F0_14_12 ( .D(\din[12][14] ), .G(n38), .Q(\q[12][14] ) );
    LD1 F0_0_12 ( .D(\din[12][0] ), .G(n38), .Q(\q[12][0] ) );
    LD1 F0_12_0 ( .D(\din[0][12] ), .G(n38), .Q(\q[0][12] ) );
    LD1 F0_2_8 ( .D(\din[8][2] ), .G(n38), .Q(\q[8][2] ) );
    LD1 F0_0_4 ( .D(\din[4][0] ), .G(n38), .Q(\q[4][0] ) );
    LD1 F0_0_3 ( .D(\din[3][0] ), .G(n38), .Q(\q[3][0] ) );
    LD1 F0_13_0 ( .D(\din[0][13] ), .G(n38), .Q(\q[0][13] ) );
    LD1 F0_4_2 ( .D(\din[2][4] ), .G(n38), .Q(\q[2][4] ) );
    LD1 F0_3_8 ( .D(\din[8][3] ), .G(n38), .Q(\q[8][3] ) );
    LD1 F0_9_5 ( .D(\din[5][9] ), .G(n38), .Q(\q[5][9] ) );
    LD1 F0_1_13 ( .D(\din[13][1] ), .G(n38), .Q(\q[13][1] ) );
    LD1 F0_1_4 ( .D(\din[4][1] ), .G(n38), .Q(\q[4][1] ) );
    LD1 F0_15_13 ( .D(\din[13][15] ), .G(n38), .Q(\q[13][15] ) );
    LD1 F0_5_10 ( .D(\din[10][5] ), .G(n38), .Q(\q[10][5] ) );
    LD1 F0_11_10 ( .D(\din[10][11] ), .G(n38), .Q(\q[10][11] ) );
    LD1 F0_6_5 ( .D(\din[5][6] ), .G(n38), .Q(\q[5][6] ) );
    LD1 F0_3_15 ( .D(\din[15][3] ), .G(n38), .Q(\q[15][3] ) );
    LD1 F0_3_3 ( .D(\din[3][3] ), .G(n38), .Q(\q[3][3] ) );
    LD1 F0_11_7 ( .D(\din[7][11] ), .G(n38), .Q(\q[7][11] ) );
    LD1 F0_9_13 ( .D(\din[13][9] ), .G(n38), .Q(\q[13][9] ) );
    LD1 F0_14_1 ( .D(\din[1][14] ), .G(n38), .Q(\q[1][14] ) );
    LD1 F0_4_9 ( .D(\din[9][4] ), .G(n38), .Q(\q[9][4] ) );
    LD1 F0_4_11 ( .D(\din[11][4] ), .G(n38), .Q(\q[11][4] ) );
    LD1 F0_10_11 ( .D(\din[11][10] ), .G(n38), .Q(\q[11][10] ) );
    LD1 F0_7_5 ( .D(\din[5][7] ), .G(n38), .Q(\q[5][7] ) );
    LD1 F0_15_1 ( .D(\din[1][15] ), .G(n38), .Q(\q[1][15] ) );
    LD1 F0_10_7 ( .D(\din[7][10] ), .G(n38), .Q(\q[7][10] ) );
    LD1 F0_5_9 ( .D(\din[9][5] ), .G(n38), .Q(\q[9][5] ) );
    LD1 F0_2_3 ( .D(\din[3][2] ), .G(n38), .Q(\q[3][2] ) );
    LD1 F0_8_12 ( .D(\din[12][8] ), .G(n38), .Q(\q[12][8] ) );
    LD1 F0_2_14 ( .D(\din[14][2] ), .G(n38), .Q(\q[14][2] ) );
    LD1 F0_15_11 ( .D(\din[11][15] ), .G(n38), .Q(\q[11][15] ) );
    LD1 F0_13_2 ( .D(\din[2][13] ), .G(n38), .Q(\q[2][13] ) );
    LD1 F0_9_7 ( .D(\din[7][9] ), .G(n38), .Q(\q[7][9] ) );
    LD1 F0_14_8 ( .D(\din[8][14] ), .G(n38), .Q(\q[8][14] ) );
    LD1 F0_13_14 ( .D(\din[14][13] ), .G(n38), .Q(\q[14][13] ) );
    LD1 F0_4_0 ( .D(\din[0][4] ), .G(n38), .Q(\q[0][4] ) );
    LD1 F0_1_11 ( .D(\din[11][1] ), .G(n38), .Q(\q[11][1] ) );
    LD1 F0_0_2 ( .D(\din[2][0] ), .G(n38), .Q(\q[2][0] ) );
    LD1 F0_7_14 ( .D(\din[14][7] ), .G(n38), .Q(\q[14][7] ) );
    LD1 F0_12_2 ( .D(\din[2][12] ), .G(n38), .Q(\q[2][12] ) );
    LD1 F0_1_6 ( .D(\din[6][1] ), .G(n38), .Q(\q[6][1] ) );
    LD1 F0_14_10 ( .D(\din[10][14] ), .G(n38), .Q(\q[10][14] ) );
    LD1 F0_5_0 ( .D(\din[0][5] ), .G(n38), .Q(\q[0][5] ) );
    LD1 F0_15_8 ( .D(\din[8][15] ), .G(n38), .Q(\q[8][15] ) );
    LD1 F0_12_15 ( .D(\din[15][12] ), .G(n38), .Q(\q[15][12] ) );
    LD1 F0_8_7 ( .D(\din[7][8] ), .G(n38), .Q(\q[7][8] ) );
    LD1 F0_6_15 ( .D(\din[15][6] ), .G(n38), .Q(\q[15][6] ) );
    LD1 F0_12_12 ( .D(\din[12][12] ), .G(n38), .Q(\q[12][12] ) );
    LD1 F0_12_5 ( .D(\din[5][12] ), .G(n38), .Q(\q[5][12] ) );
    LD1 F0_8_0 ( .D(\din[0][8] ), .G(n38), .Q(\q[0][8] ) );
    LD1 F0_6_12 ( .D(\din[12][6] ), .G(n38), .Q(\q[12][6] ) );
    LD1 F0_10_9 ( .D(\din[9][10] ), .G(n38), .Q(\q[9][10] ) );
    LD1 F0_5_7 ( .D(\din[7][5] ), .G(n38), .Q(\q[7][5] ) );
    LD1 F0_0_10 ( .D(\din[10][0] ), .G(n38), .Q(\q[10][0] ) );
    LD1 F0_0_6 ( .D(\din[6][0] ), .G(n38), .Q(\q[6][0] ) );
    LD1 F0_13_5 ( .D(\din[5][13] ), .G(n38), .Q(\q[5][13] ) );
    LD1 F0_11_9 ( .D(\din[9][11] ), .G(n38), .Q(\q[9][11] ) );
    LD1 F0_7_13 ( .D(\din[13][7] ), .G(n38), .Q(\q[13][7] ) );
    LD1 F0_1_1 ( .D(\din[1][1] ), .G(n38), .Q(\q[1][1] ) );
    LD1 F0_13_13 ( .D(\din[13][13] ), .G(n38), .Q(\q[13][13] ) );
    LD1 F0_9_0 ( .D(\din[0][9] ), .G(n38), .Q(\q[0][9] ) );
    LD1 F0_4_7 ( .D(\din[7][4] ), .G(n38), .Q(\q[7][4] ) );
    LD1 F0_8_15 ( .D(\din[15][8] ), .G(n38), .Q(\q[15][8] ) );
    LD1 F0_8_9 ( .D(\din[9][8] ), .G(n38), .Q(\q[9][8] ) );
    LD1 F0_7_2 ( .D(\din[2][7] ), .G(n38), .Q(\q[2][7] ) );
    LD1 F0_2_13 ( .D(\din[13][2] ), .G(n38), .Q(\q[13][2] ) );
    LD1 F0_2_4 ( .D(\din[4][2] ), .G(n38), .Q(\q[4][2] ) );
    LD1 F0_10_0 ( .D(\din[0][10] ), .G(n38), .Q(\q[0][10] ) );
    LD1 F0_15_6 ( .D(\din[6][15] ), .G(n38), .Q(\q[6][15] ) );
    LD1 F0_3_4 ( .D(\din[4][3] ), .G(n38), .Q(\q[4][3] ) );
    LD1 F0_6_2 ( .D(\din[2][6] ), .G(n38), .Q(\q[2][6] ) );
    LD1 F0_14_6 ( .D(\din[6][14] ), .G(n38), .Q(\q[6][14] ) );
    LD1 F0_11_0 ( .D(\din[0][11] ), .G(n38), .Q(\q[0][11] ) );
    LD1 F0_9_14 ( .D(\din[14][9] ), .G(n38), .Q(\q[14][9] ) );
    LD1 F0_3_12 ( .D(\din[12][3] ), .G(n38), .Q(\q[12][3] ) );
    LD1 F0_9_9 ( .D(\din[9][9] ), .G(n38), .Q(\q[9][9] ) );
    LD1 F0_9_1 ( .D(\din[1][9] ), .G(n38), .Q(\q[1][9] ) );
    LD1 F0_13_4 ( .D(\din[4][13] ), .G(n38), .Q(\q[4][13] ) );
    LD1 F0_1_8 ( .D(\din[8][1] ), .G(n38), .Q(\q[8][1] ) );
    LD1 F0_1_0 ( .D(\din[0][1] ), .G(n38), .Q(\q[0][1] ) );
    LD1 F0_0_8 ( .D(\din[8][0] ), .G(n38), .Q(\q[8][0] ) );
    LD1 F0_11_8 ( .D(\din[8][11] ), .G(n38), .Q(\q[8][11] ) );
    LD1 F0_13_12 ( .D(\din[12][13] ), .G(n38), .Q(\q[12][13] ) );
    LD1 F0_7_12 ( .D(\din[12][7] ), .G(n38), .Q(\q[12][7] ) );
    LD1 F0_12_4 ( .D(\din[4][12] ), .G(n38), .Q(\q[4][12] ) );
    LD1 F0_4_6 ( .D(\din[6][4] ), .G(n38), .Q(\q[6][4] ) );
    LD1 F0_5_6 ( .D(\din[6][5] ), .G(n38), .Q(\q[6][5] ) );
    LD1 F0_10_8 ( .D(\din[8][10] ), .G(n38), .Q(\q[8][10] ) );
    LD1 F0_0_1 ( .D(\din[1][0] ), .G(n38), .Q(\q[1][0] ) );
    LD1 F0_12_13 ( .D(\din[13][12] ), .G(n38), .Q(\q[13][12] ) );
    LD1 F0_9_8 ( .D(\din[8][9] ), .G(n38), .Q(\q[8][9] ) );
    LD1 F0_8_1 ( .D(\din[1][8] ), .G(n38), .Q(\q[1][8] ) );
    LD1 F0_6_13 ( .D(\din[13][6] ), .G(n38), .Q(\q[13][6] ) );
    LD1 F0_6_3 ( .D(\din[3][6] ), .G(n38), .Q(\q[3][6] ) );
    LD1 F0_14_7 ( .D(\din[7][14] ), .G(n38), .Q(\q[7][14] ) );
    LD1 F0_11_1 ( .D(\din[1][11] ), .G(n38), .Q(\q[1][11] ) );
    LD1 F0_9_15 ( .D(\din[15][9] ), .G(n38), .Q(\q[15][9] ) );
    LD1 F0_3_13 ( .D(\din[13][3] ), .G(n38), .Q(\q[13][3] ) );
    LD1 F0_3_5 ( .D(\din[5][3] ), .G(n38), .Q(\q[5][3] ) );
    LD1 F0_7_3 ( .D(\din[3][7] ), .G(n38), .Q(\q[3][7] ) );
    LD1 F0_2_5 ( .D(\din[5][2] ), .G(n38), .Q(\q[5][2] ) );
    LD1 F0_1_9 ( .D(\din[9][1] ), .G(n38), .Q(\q[9][1] ) );
    LD1 F0_15_7 ( .D(\din[7][15] ), .G(n38), .Q(\q[7][15] ) );
    LD1 F0_10_1 ( .D(\din[1][10] ), .G(n38), .Q(\q[1][10] ) );
    LD1 F0_8_14 ( .D(\din[14][8] ), .G(n38), .Q(\q[14][8] ) );
    LD1 F0_8_8 ( .D(\din[8][8] ), .G(n38), .Q(\q[8][8] ) );
    LD1 F0_8_13 ( .D(\din[13][8] ), .G(n38), .Q(\q[13][8] ) );
    LD1 F0_4_10 ( .D(\din[10][4] ), .G(n38), .Q(\q[10][4] ) );
    LD1 F0_2_15 ( .D(\din[15][2] ), .G(n38), .Q(\q[15][2] ) );
    LD1 F0_2_12 ( .D(\din[12][2] ), .G(n38), .Q(\q[12][2] ) );
    LD1 F0_10_10 ( .D(\din[10][10] ), .G(n38), .Q(\q[10][10] ) );
    LD1 F0_15_0 ( .D(\din[0][15] ), .G(n38), .Q(\q[0][15] ) );
    LD1 F0_7_4 ( .D(\din[4][7] ), .G(n38), .Q(\q[4][7] ) );
    LD1 F0_5_8 ( .D(\din[8][5] ), .G(n38), .Q(\q[8][5] ) );
    LD1 F0_2_2 ( .D(\din[2][2] ), .G(n38), .Q(\q[2][2] ) );
    LD1 F0_10_6 ( .D(\din[6][10] ), .G(n38), .Q(\q[6][10] ) );
    LD1 F0_6_4 ( .D(\din[4][6] ), .G(n38), .Q(\q[4][6] ) );
    LD1 F0_3_14 ( .D(\din[14][3] ), .G(n38), .Q(\q[14][3] ) );
    LD1 F0_3_2 ( .D(\din[2][3] ), .G(n38), .Q(\q[2][3] ) );
    LD1 F0_0_9 ( .D(\din[9][0] ), .G(n38), .Q(\q[9][0] ) );
    LD1 F0_11_6 ( .D(\din[6][11] ), .G(n38), .Q(\q[6][11] ) );
    LD1 F0_14_0 ( .D(\din[0][14] ), .G(n38), .Q(\q[0][14] ) );
    LD1 F0_9_12 ( .D(\din[12][9] ), .G(n38), .Q(\q[12][9] ) );
    LD1 F0_5_11 ( .D(\din[11][5] ), .G(n38), .Q(\q[11][5] ) );
    LD1 F0_11_11 ( .D(\din[11][11] ), .G(n38), .Q(\q[11][11] ) );
    LD1 F0_12_14 ( .D(\din[14][12] ), .G(n38), .Q(\q[14][12] ) );
    LD1 F0_8_6 ( .D(\din[6][8] ), .G(n38), .Q(\q[6][8] ) );
    LD1 F0_14_11 ( .D(\din[11][14] ), .G(n38), .Q(\q[11][14] ) );
    LD1 F0_12_3 ( .D(\din[3][12] ), .G(n38), .Q(\q[3][12] ) );
    LD1 F0_6_14 ( .D(\din[14][6] ), .G(n38), .Q(\q[14][6] ) );
    LD1 F0_4_8 ( .D(\din[8][4] ), .G(n38), .Q(\q[8][4] ) );
    LD1 F0_15_9 ( .D(\din[9][15] ), .G(n38), .Q(\q[9][15] ) );
    LD1 F0_5_1 ( .D(\din[1][5] ), .G(n38), .Q(\q[1][5] ) );
    LD1 F0_14_9 ( .D(\din[9][14] ), .G(n38), .Q(\q[9][14] ) );
    LD1 F0_13_3 ( .D(\din[3][13] ), .G(n38), .Q(\q[3][13] ) );
    LD1 F0_13_15 ( .D(\din[15][13] ), .G(n38), .Q(\q[15][13] ) );
    LD1 F0_7_15 ( .D(\din[15][7] ), .G(n38), .Q(\q[15][7] ) );
    LD1 F0_4_1 ( .D(\din[1][4] ), .G(n38), .Q(\q[1][4] ) );
    LD1 F0_0_11 ( .D(\din[11][0] ), .G(n38), .Q(\q[11][0] ) );
    LD1 F0_0_7 ( .D(\din[7][0] ), .G(n38), .Q(\q[7][0] ) );
    LD1 F0_0_0 ( .D(\din[0][0] ), .G(n38), .Q(\q[0][0] ) );
    LD1 F0_1_7 ( .D(\din[7][1] ), .G(n38), .Q(\q[7][1] ) );
    LD1 F0_15_10 ( .D(\din[10][15] ), .G(n38), .Q(\q[10][15] ) );
    LD1 F0_9_6 ( .D(\din[6][9] ), .G(n38), .Q(\q[6][9] ) );
    LD1 F0_1_10 ( .D(\din[10][1] ), .G(n38), .Q(\q[10][1] ) );
    NR2 U72 ( .A(n60), .B(wr_n), .Z(\wren[6] ) );
    NR2 U73 ( .A(n61), .B(wr_n), .Z(\wren[1] ) );
    NR2 U74 ( .A(n62), .B(wr_n), .Z(\wren[8] ) );
    NR2 U75 ( .A(n63), .B(wr_n), .Z(\wren[10] ) );
    NR2 U76 ( .A(n64), .B(wr_n), .Z(\wren[0] ) );
    NR2 U77 ( .A(n65), .B(wr_n), .Z(\wren[11] ) );
    NR2 U78 ( .A(n66), .B(wr_n), .Z(\wren[9] ) );
    NR2 U79 ( .A(n67), .B(wr_n), .Z(\wren[7] ) );
    NR2 U80 ( .A(n68), .B(wr_n), .Z(\wren[14] ) );
    NR2 U81 ( .A(n69), .B(wr_n), .Z(\wren[5] ) );
    NR2 U82 ( .A(n70), .B(wr_n), .Z(\wren[2] ) );
    NR2 U83 ( .A(n71), .B(wr_n), .Z(\wren[13] ) );
    NR2 U84 ( .A(n72), .B(wr_n), .Z(\wren[3] ) );
    NR2 U85 ( .A(n73), .B(wr_n), .Z(\wren[12] ) );
    NR2 U86 ( .A(n108), .B(wr_n), .Z(\wren[15] ) );
    NR2 U87 ( .A(n109), .B(wr_n), .Z(\wren[4] ) );
    IV U88 ( .A(clk), .Z(n38) );
    IV U89 ( .A(wr_addr[9]), .Z(n66) );
    IV U90 ( .A(wr_addr[8]), .Z(n62) );
    IV U91 ( .A(wr_addr[7]), .Z(n67) );
    IV U92 ( .A(wr_addr[6]), .Z(n60) );
    IV U93 ( .A(wr_addr[5]), .Z(n69) );
    IV U94 ( .A(wr_addr[4]), .Z(n109) );
    IV U95 ( .A(wr_addr[3]), .Z(n72) );
    IV U96 ( .A(wr_addr[2]), .Z(n70) );
    IV U97 ( .A(wr_addr[1]), .Z(n61) );
    IV U98 ( .A(wr_addr[15]), .Z(n108) );
    IV U99 ( .A(wr_addr[14]), .Z(n68) );
    IV U100 ( .A(wr_addr[13]), .Z(n71) );
    IV U101 ( .A(wr_addr[12]), .Z(n73) );
    IV U102 ( .A(wr_addr[11]), .Z(n65) );
    IV U103 ( .A(wr_addr[10]), .Z(n63) );
    IV U104 ( .A(wr_addr[0]), .Z(n64) );
endmodule


module fifo_DW01_mux_any_256_4_16_0 ( A, SEL, MUX );
input  [255:0] A;
input  [3:0] SEL;
output [15:0] MUX;
    wire \tmp[3][136] , \tmp[3][14] , \tmp[3][132] , \tmp[3][10] , 
        \tmp[3][139] , \tmp[3][130] , \tmp[3][129] , \tmp[3][12] , 
        \tmp[3][134] , \tmp[3][1] , \tmp[3][8] , \tmp[3][141] , \tmp[3][5] , 
        \tmp[3][7] , \tmp[3][143] , \tmp[3][3] , \tmp[3][142] , \tmp[3][2] , 
        \tmp[3][6] , \tmp[3][4] , \tmp[3][0] , \tmp[3][9] , \tmp[3][140] , 
        \tmp[3][135] , \tmp[3][138] , \tmp[3][13] , \tmp[3][131] , 
        \tmp[3][128] , \tmp[3][11] , \tmp[3][133] , \tmp[3][137] , 
        \tmp[3][15] , n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
        n85, n86, n87, n88, n89, n90;
    MUX81P MX8_1_1_0 ( .D0(A[0]), .D1(A[16]), .D2(A[32]), .D3(A[48]), .D4(A
        [64]), .D5(A[80]), .D6(A[96]), .D7(A[112]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][0] ) );
    MUX81P MX8_1_1_1 ( .D0(A[1]), .D1(A[17]), .D2(A[33]), .D3(A[49]), .D4(A
        [65]), .D5(A[81]), .D6(A[97]), .D7(A[113]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][1] ) );
    MUX81P MX8_1_1_2 ( .D0(A[2]), .D1(A[18]), .D2(A[34]), .D3(A[50]), .D4(A
        [66]), .D5(A[82]), .D6(A[98]), .D7(A[114]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][2] ) );
    MUX81P MX8_1_5_10 ( .D0(A[138]), .D1(A[154]), .D2(A[170]), .D3(A[186]), 
        .D4(A[202]), .D5(A[218]), .D6(A[234]), .D7(A[250]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][138] ) );
    MUX81P MX8_1_1_3 ( .D0(A[3]), .D1(A[19]), .D2(A[35]), .D3(A[51]), .D4(A
        [67]), .D5(A[83]), .D6(A[99]), .D7(A[115]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][3] ) );
    MUX81P MX8_1_1_4 ( .D0(A[4]), .D1(A[20]), .D2(A[36]), .D3(A[52]), .D4(A
        [68]), .D5(A[84]), .D6(A[100]), .D7(A[116]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][4] ) );
    MUX81P MX8_1_1_5 ( .D0(A[5]), .D1(A[21]), .D2(A[37]), .D3(A[53]), .D4(A
        [69]), .D5(A[85]), .D6(A[101]), .D7(A[117]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][5] ) );
    MUX81P MX8_1_1_11 ( .D0(A[11]), .D1(A[27]), .D2(A[43]), .D3(A[59]), .D4(A
        [75]), .D5(A[91]), .D6(A[107]), .D7(A[123]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][11] ) );
    MUX81P MX8_1_5_3 ( .D0(A[131]), .D1(A[147]), .D2(A[163]), .D3(A[179]), 
        .D4(A[195]), .D5(A[211]), .D6(A[227]), .D7(A[243]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][131] ) );
    MUX81P MX8_1_5_4 ( .D0(A[132]), .D1(A[148]), .D2(A[164]), .D3(A[180]), 
        .D4(A[196]), .D5(A[212]), .D6(A[228]), .D7(A[244]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][132] ) );
    MUX81P MX8_1_1_10 ( .D0(A[10]), .D1(A[26]), .D2(A[42]), .D3(A[58]), .D4(A
        [74]), .D5(A[90]), .D6(A[106]), .D7(A[122]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][10] ) );
    MUX81P MX8_1_5_2 ( .D0(A[130]), .D1(A[146]), .D2(A[162]), .D3(A[178]), 
        .D4(A[194]), .D5(A[210]), .D6(A[226]), .D7(A[242]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][130] ) );
    MUX81P MX8_1_5_5 ( .D0(A[133]), .D1(A[149]), .D2(A[165]), .D3(A[181]), 
        .D4(A[197]), .D5(A[213]), .D6(A[229]), .D7(A[245]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][133] ) );
    MUX81P MX8_1_5_11 ( .D0(A[139]), .D1(A[155]), .D2(A[171]), .D3(A[187]), 
        .D4(A[203]), .D5(A[219]), .D6(A[235]), .D7(A[251]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][139] ) );
    MUX81P MX8_1_1_8 ( .D0(A[8]), .D1(A[24]), .D2(A[40]), .D3(A[56]), .D4(A
        [72]), .D5(A[88]), .D6(A[104]), .D7(A[120]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][8] ) );
    MUX81P MX8_1_5_13 ( .D0(A[141]), .D1(A[157]), .D2(A[173]), .D3(A[189]), 
        .D4(A[205]), .D5(A[221]), .D6(A[237]), .D7(A[253]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][141] ) );
    MUX81P MX8_1_1_6 ( .D0(A[6]), .D1(A[22]), .D2(A[38]), .D3(A[54]), .D4(A
        [70]), .D5(A[86]), .D6(A[102]), .D7(A[118]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][6] ) );
    MUX81P MX8_1_1_12 ( .D0(A[12]), .D1(A[28]), .D2(A[44]), .D3(A[60]), .D4(A
        [76]), .D5(A[92]), .D6(A[108]), .D7(A[124]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][12] ) );
    MUX81P MX8_1_1_15 ( .D0(A[15]), .D1(A[31]), .D2(A[47]), .D3(A[63]), .D4(A
        [79]), .D5(A[95]), .D6(A[111]), .D7(A[127]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][15] ) );
    MUX81P MX8_1_5_0 ( .D0(A[128]), .D1(A[144]), .D2(A[160]), .D3(A[176]), 
        .D4(A[192]), .D5(A[208]), .D6(A[224]), .D7(A[240]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][128] ) );
    MUX81P MX8_1_5_7 ( .D0(A[135]), .D1(A[151]), .D2(A[167]), .D3(A[183]), 
        .D4(A[199]), .D5(A[215]), .D6(A[231]), .D7(A[247]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][135] ) );
    MUX81P MX8_1_1_7 ( .D0(A[7]), .D1(A[23]), .D2(A[39]), .D3(A[55]), .D4(A
        [71]), .D5(A[87]), .D6(A[103]), .D7(A[119]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][7] ) );
    MUX81P MX8_1_5_9 ( .D0(A[137]), .D1(A[153]), .D2(A[169]), .D3(A[185]), 
        .D4(A[201]), .D5(A[217]), .D6(A[233]), .D7(A[249]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][137] ) );
    MUX81P MX8_1_5_14 ( .D0(A[142]), .D1(A[158]), .D2(A[174]), .D3(A[190]), 
        .D4(A[206]), .D5(A[222]), .D6(A[238]), .D7(A[254]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][142] ) );
    MUX81P MX8_1_1_9 ( .D0(A[9]), .D1(A[25]), .D2(A[41]), .D3(A[57]), .D4(A
        [73]), .D5(A[89]), .D6(A[105]), .D7(A[121]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][9] ) );
    MUX81P MX8_1_1_14 ( .D0(A[14]), .D1(A[30]), .D2(A[46]), .D3(A[62]), .D4(A
        [78]), .D5(A[94]), .D6(A[110]), .D7(A[126]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][14] ) );
    MUX81P MX8_1_5_1 ( .D0(A[129]), .D1(A[145]), .D2(A[161]), .D3(A[177]), 
        .D4(A[193]), .D5(A[209]), .D6(A[225]), .D7(A[241]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][129] ) );
    MUX81P MX8_1_5_8 ( .D0(A[136]), .D1(A[152]), .D2(A[168]), .D3(A[184]), 
        .D4(A[200]), .D5(A[216]), .D6(A[232]), .D7(A[248]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][136] ) );
    MUX81P MX8_1_5_15 ( .D0(A[143]), .D1(A[159]), .D2(A[175]), .D3(A[191]), 
        .D4(A[207]), .D5(A[223]), .D6(A[239]), .D7(A[255]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][143] ) );
    MUX81P MX8_1_5_12 ( .D0(A[140]), .D1(A[156]), .D2(A[172]), .D3(A[188]), 
        .D4(A[204]), .D5(A[220]), .D6(A[236]), .D7(A[252]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][140] ) );
    MUX81P MX8_1_1_13 ( .D0(A[13]), .D1(A[29]), .D2(A[45]), .D3(A[61]), .D4(A
        [77]), .D5(A[93]), .D6(A[109]), .D7(A[125]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][13] ) );
    MUX81P MX8_1_5_6 ( .D0(A[134]), .D1(A[150]), .D2(A[166]), .D3(A[182]), 
        .D4(A[198]), .D5(A[214]), .D6(A[230]), .D7(A[246]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][134] ) );
    AO2 U72 ( .A(\tmp[3][9] ), .B(n75), .C(\tmp[3][137] ), .D(SEL[3]), .Z(n74)
         );
    AO2 U73 ( .A(\tmp[3][8] ), .B(n75), .C(\tmp[3][136] ), .D(SEL[3]), .Z(n76)
         );
    AO2 U74 ( .A(\tmp[3][7] ), .B(n75), .C(\tmp[3][135] ), .D(SEL[3]), .Z(n77)
         );
    AO2 U75 ( .A(\tmp[3][6] ), .B(n75), .C(\tmp[3][134] ), .D(SEL[3]), .Z(n78)
         );
    AO2 U76 ( .A(\tmp[3][5] ), .B(n75), .C(\tmp[3][133] ), .D(SEL[3]), .Z(n79)
         );
    AO2 U77 ( .A(\tmp[3][4] ), .B(n75), .C(\tmp[3][132] ), .D(SEL[3]), .Z(n80)
         );
    AO2 U78 ( .A(\tmp[3][3] ), .B(n75), .C(\tmp[3][131] ), .D(SEL[3]), .Z(n81)
         );
    AO2 U79 ( .A(\tmp[3][2] ), .B(n75), .C(\tmp[3][130] ), .D(SEL[3]), .Z(n82)
         );
    AO2 U80 ( .A(\tmp[3][1] ), .B(n75), .C(\tmp[3][129] ), .D(SEL[3]), .Z(n83)
         );
    AO2 U81 ( .A(\tmp[3][15] ), .B(n75), .C(\tmp[3][143] ), .D(SEL[3]), .Z(n84
        ) );
    AO2 U82 ( .A(\tmp[3][14] ), .B(n75), .C(\tmp[3][142] ), .D(SEL[3]), .Z(n85
        ) );
    AO2 U83 ( .A(\tmp[3][13] ), .B(n75), .C(\tmp[3][141] ), .D(SEL[3]), .Z(n86
        ) );
    AO2 U84 ( .A(\tmp[3][12] ), .B(n75), .C(\tmp[3][140] ), .D(SEL[3]), .Z(n87
        ) );
    AO2 U85 ( .A(\tmp[3][11] ), .B(n75), .C(\tmp[3][139] ), .D(SEL[3]), .Z(n88
        ) );
    AO2 U86 ( .A(\tmp[3][10] ), .B(n75), .C(\tmp[3][138] ), .D(SEL[3]), .Z(n89
        ) );
    AO2 U87 ( .A(\tmp[3][0] ), .B(n75), .C(\tmp[3][128] ), .D(SEL[3]), .Z(n90)
         );
    IV U88 ( .A(SEL[3]), .Z(n75) );
    IV U89 ( .A(n74), .Z(MUX[9]) );
    IV U90 ( .A(n76), .Z(MUX[8]) );
    IV U91 ( .A(n77), .Z(MUX[7]) );
    IV U92 ( .A(n78), .Z(MUX[6]) );
    IV U93 ( .A(n79), .Z(MUX[5]) );
    IV U94 ( .A(n80), .Z(MUX[4]) );
    IV U95 ( .A(n81), .Z(MUX[3]) );
    IV U96 ( .A(n82), .Z(MUX[2]) );
    IV U97 ( .A(n83), .Z(MUX[1]) );
    IV U98 ( .A(n84), .Z(MUX[15]) );
    IV U99 ( .A(n85), .Z(MUX[14]) );
    IV U100 ( .A(n86), .Z(MUX[13]) );
    IV U101 ( .A(n87), .Z(MUX[12]) );
    IV U102 ( .A(n88), .Z(MUX[11]) );
    IV U103 ( .A(n89), .Z(MUX[10]) );
    IV U104 ( .A(n90), .Z(MUX[0]) );
endmodule


module fifo_DW_MEM_R_W_S_LAT_16_16_0 ( clk, wr_n, rd_addr, wr_addr, data_in, 
    data_out );
output [15:0] data_out;
input  [3:0] rd_addr;
input  [15:0] wr_addr;
input  [15:0] data_in;
input  clk, wr_n;
    wire \q[15][15] , \q[15][14] , \q[15][12] , \q[15][9] , \q[15][6] , 
        \q[15][2] , \q[14][1] , \q[10][15] , \q[6][0] , \q[1][12] , 
        \din[15][0] , \q[11][13] , \q[11][9] , \q[10][3] , \din[11][2] , 
        \din[5][1] , \din[1][3] , \q[2][2] , \din[6][12] , \q[9][14] , 
        \q[8][4] , \din[0][9] , \din[10][8] , \q[6][10] , \q[3][8] , \q[3][1] , 
        \din[10][10] , \din[8][10] , \q[0][14] , \q[11][0] , \din[10][1] , 
        \din[14][3] , \din[0][0] , \din[4][2] , \q[14][8] , \q[7][3] , 
        \din[7][14] , \din[1][10] , \q[14][5] , \q[10][7] , \q[9][10] , 
        \q[9][7] , \q[8][12] , \q[6][9] , \din[15][9] , \din[5][8] , \q[8][0] , 
        \din[10][14] , \din[8][14] , \q[2][6] , \din[11][6] , \din[0][12] , 
        \din[15][4] , \din[1][7] , \din[5][5] , \q[10][11] , \q[7][12] , 
        \q[9][3] , \q[6][4] , \din[9][12] , \q[7][7] , \din[11][12] , 
        \din[14][7] , \din[7][10] , \din[1][14] , \q[15][4] , \q[11][4] , 
        \q[8][9] , \din[10][5] , \din[4][6] , \din[0][4] , \q[7][5] , 
        \q[6][14] , \q[3][5] , \q[0][10] , \din[14][5] , \din[7][12] , 
        \din[4][4] , \q[15][0] , \q[14][7] , \q[11][15] , \q[11][6] , 
        \din[10][7] , \q[3][7] , \din[0][6] , \q[0][12] , \q[10][5] , 
        \q[9][8] , \q[9][1] , \q[8][14] , \din[11][10] , \din[9][10] , 
        \q[2][4] , \din[6][14] , \din[0][10] , \din[11][4] , \din[1][5] , 
        \din[15][6] , \q[11][11] , \q[10][13] , \q[6][6] , \din[5][7] , 
        \q[10][8] , \q[9][12] , \q[8][2] , \q[7][10] , \q[1][14] , \q[8][10] , 
        \q[2][9] , \din[11][14] , \din[9][14] , \q[9][5] , \din[1][8] , 
        \q[3][3] , \din[11][9] , \q[11][2] , \q[6][12] , \din[10][3] , 
        \din[0][2] , \din[14][1] , \q[8][6] , \q[7][1] , \din[4][0] , 
        \din[1][12] , \q[7][8] , \din[10][12] , \q[14][3] , \q[7][14] , 
        \q[1][10] , \din[14][8] , \din[8][12] , \din[4][9] , \q[6][2] , 
        \din[15][2] , \din[5][3] , \q[12][7] , \q[10][1] , \din[11][0] , 
        \q[4][4] , \q[2][0] , \din[1][1] , \wren[8] , \din[6][10] , 
        \din[0][14] , \din[5][11] , \din[3][15] , \din[7][5] , \q[0][6] , 
        \din[13][6] , \din[3][7] , \q[14][14] , \q[13][4] , \q[4][15] , 
        \q[2][11] , \q[1][5] , \din[13][13] , \din[9][1] , \din[2][13] , 
        \din[9][8] , \din[2][4] , \q[12][10] , \q[5][13] , \din[12][5] , 
        \din[6][6] , \q[14][12] , \q[14][10] , \q[13][12] , \q[13][9] , 
        \q[5][7] , \q[1][8] , \wren[1] , \din[14][11] , \din[12][15] , 
        \din[15][13] , \din[8][2] , \din[12][8] , \din[9][5] , \q[4][11] , 
        \q[2][15] , \din[2][9] , \q[12][3] , \q[0][2] , \din[3][3] , \q[4][9] , 
        \q[4][0] , \din[13][2] , \din[7][1] , \din[8][6] , \din[5][15] , 
        \din[3][11] , \wren[5] , \din[14][15] , \din[12][11] , \din[7][8] , 
        \q[13][0] , \q[12][14] , \q[5][3] , \q[3][13] , \din[6][2] , 
        \q[5][15] , \q[1][1] , \wren[13] , \din[2][0] , \din[12][1] , 
        \din[4][13] , \q[3][11] , \q[13][10] , \q[13][2] , \q[5][1] , 
        \wren[11] , \din[6][0] , \din[2][2] , \q[12][8] , \q[1][3] , 
        \din[12][3] , \din[4][11] , \din[2][15] , \din[13][9] , \q[0][9] , 
        \din[3][8] , \q[0][0] , \wren[7] , \din[12][13] , \din[8][4] , 
        \q[15][11] , \q[15][10] , \q[13][6] , \q[12][1] , \q[4][13] , 
        \q[5][8] , \q[4][2] , \din[13][0] , \din[3][1] , \din[7][3] , 
        \din[3][13] , \din[6][9] , \q[1][7] , \wren[3] , \din[15][11] , 
        \din[9][7] , \din[13][15] , \din[14][13] , \din[8][0] , \din[4][15] , 
        \din[2][11] , \q[12][12] , \wren[15] , \din[2][6] , \din[12][7] , 
        \din[6][4] , \q[12][5] , \q[5][11] , \q[3][15] , \q[5][5] , \q[4][6] , 
        \din[15][15] , \din[13][11] , \din[9][3] , \din[7][7] , \din[5][13] , 
        \din[3][5] , \q[2][13] , \din[13][4] , \q[13][15] , \q[13][14] , 
        \q[13][7] , \q[0][4] , \wren[14] , \wren[2] , \din[8][9] , 
        \din[14][12] , \din[8][1] , \q[12][13] , \q[1][6] , \din[12][6] , 
        \din[2][7] , \din[4][14] , \din[2][10] , \q[5][10] , \q[5][4] , 
        \q[3][14] , \q[4][7] , \din[15][14] , \din[6][5] , \din[13][10] , 
        \din[9][2] , \din[7][6] , \din[5][12] , \q[2][12] , \q[0][5] , 
        \din[8][8] , \q[14][13] , \q[12][4] , \din[3][4] , \q[5][14] , 
        \q[3][10] , \din[13][5] , \din[6][1] , \q[13][3] , \q[5][0] , 
        \q[1][2] , \din[4][10] , \din[2][14] , \din[2][3] , \q[12][9] , 
        \q[0][8] , \wren[10] , \din[12][2] , \din[8][5] , \din[13][8] , 
        \q[12][0] , \wren[6] , \din[12][12] , \din[3][9] , \din[13][1] , 
        \din[3][0] , \q[15][13] , \q[14][11] , \q[13][13] , \q[13][11] , 
        \q[13][8] , \q[5][9] , \q[4][12] , \q[4][3] , \q[0][1] , \din[7][2] , 
        \din[3][12] , \din[15][10] , \din[13][14] , \din[9][6] , \din[6][8] , 
        \din[12][9] , \q[12][2] , \q[1][9] , \din[15][12] , \din[2][8] , 
        \din[9][4] , \din[3][2] , \q[4][10] , \q[0][3] , \din[13][3] , 
        \q[2][14] , \q[12][15] , \q[4][8] , \q[4][1] , \din[5][14] , 
        \din[3][10] , \din[8][7] , \din[7][0] , \din[7][9] , \wren[4] , 
        \din[14][14] , \din[12][10] , \din[6][3] , \q[13][1] , \q[5][2] , 
        \q[3][12] , \q[1][0] , \din[4][12] , \wren[12] , \q[4][5] , \wren[9] , 
        \din[12][0] , \din[2][1] , \din[7][4] , \din[5][10] , \din[3][14] , 
        \q[15][8] , \q[15][1] , \q[14][15] , \q[13][5] , \q[12][6] , 
        \q[4][14] , \q[2][10] , \q[0][7] , \din[13][12] , \din[13][7] , 
        \din[3][6] , \din[9][0] , \din[2][5] , \q[5][12] , \q[1][4] , 
        \din[12][4] , \din[9][9] , \din[2][12] , \q[12][11] , \q[11][10] , 
        \q[11][3] , \q[10][9] , \q[8][11] , \q[5][6] , \din[6][7] , \wren[0] , 
        \din[14][10] , \din[12][14] , \din[8][3] , \q[9][4] , \din[9][15] , 
        \q[2][8] , \din[11][15] , \din[11][8] , \din[1][9] , \din[10][2] , 
        \din[0][3] , \q[3][2] , \q[7][0] , \q[6][13] , \din[14][0] , 
        \din[1][13] , \q[8][7] , \din[4][1] , \q[15][7] , \q[15][5] , 
        \q[14][2] , \q[7][9] , \din[14][9] , \din[8][13] , \din[4][8] , 
        \din[10][13] , \din[15][3] , \din[5][2] , \q[10][0] , \q[7][15] , 
        \q[6][3] , \q[2][1] , \q[1][11] , \din[6][11] , \din[0][15] , 
        \din[11][1] , \din[14][4] , \din[1][0] , \din[4][5] , \q[14][6] , 
        \q[11][14] , \q[7][4] , \q[3][6] , \din[7][13] , \q[0][13] , 
        \q[11][7] , \din[10][6] , \q[10][12] , \q[10][4] , \q[9][9] , 
        \q[9][0] , \din[11][11] , \din[0][7] , \q[8][15] , \din[9][11] , 
        \din[11][5] , \din[1][4] , \q[2][5] , \din[6][15] , \din[0][11] , 
        \q[7][11] , \q[1][15] , \q[6][7] , \din[15][7] , \q[14][4] , 
        \q[10][10] , \q[10][6] , \q[9][13] , \q[8][3] , \din[5][6] , 
        \q[9][11] , \q[8][1] , \din[10][15] , \din[8][15] , \din[11][7] , 
        \q[7][13] , \q[6][5] , \q[2][7] , \din[1][6] , \din[0][13] , 
        \din[15][5] , \din[5][4] , \q[9][2] , \din[11][13] , \din[9][13] , 
        \din[14][6] , \q[15][3] , \q[14][0] , \q[11][5] , \q[8][8] , \q[7][6] , 
        \din[4][7] , \q[6][15] , \q[3][4] , \din[7][11] , \din[1][15] , 
        \q[0][11] , \din[10][4] , \din[0][5] , \din[15][1] , \q[11][12] , 
        \q[11][8] , \q[10][14] , \din[5][0] , \q[10][2] , \q[6][1] , 
        \q[1][13] , \q[2][3] , \din[11][3] , \din[6][13] , \din[1][2] , 
        \q[3][9] , \q[11][1] , \q[9][15] , \q[8][5] , \din[0][8] , 
        \din[10][11] , \din[10][9] , \din[8][11] , \din[10][0] , \q[6][11] , 
        \q[3][0] , \din[0][1] , \q[0][15] , \q[7][2] , \din[14][2] , 
        \din[7][15] , \din[1][11] , \din[4][3] , \q[14][9] , \q[6][8] , 
        \q[9][6] , \q[8][13] , \din[15][8] , \din[5][9] , n73, n91, n92, n93, 
        n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107;
    fifo_DW01_mux_any_256_4_16_0 MX ( .A({\q[15][15] , \q[15][14] , 
        \q[15][13] , \q[15][12] , \q[15][11] , \q[15][10] , \q[15][9] , 
        \q[15][8] , \q[15][7] , \q[15][6] , \q[15][5] , \q[15][4] , \q[15][3] , 
        \q[15][2] , \q[15][1] , \q[15][0] , \q[14][15] , \q[14][14] , 
        \q[14][13] , \q[14][12] , \q[14][11] , \q[14][10] , \q[14][9] , 
        \q[14][8] , \q[14][7] , \q[14][6] , \q[14][5] , \q[14][4] , \q[14][3] , 
        \q[14][2] , \q[14][1] , \q[14][0] , \q[13][15] , \q[13][14] , 
        \q[13][13] , \q[13][12] , \q[13][11] , \q[13][10] , \q[13][9] , 
        \q[13][8] , \q[13][7] , \q[13][6] , \q[13][5] , \q[13][4] , \q[13][3] , 
        \q[13][2] , \q[13][1] , \q[13][0] , \q[12][15] , \q[12][14] , 
        \q[12][13] , \q[12][12] , \q[12][11] , \q[12][10] , \q[12][9] , 
        \q[12][8] , \q[12][7] , \q[12][6] , \q[12][5] , \q[12][4] , \q[12][3] , 
        \q[12][2] , \q[12][1] , \q[12][0] , \q[11][15] , \q[11][14] , 
        \q[11][13] , \q[11][12] , \q[11][11] , \q[11][10] , \q[11][9] , 
        \q[11][8] , \q[11][7] , \q[11][6] , \q[11][5] , \q[11][4] , \q[11][3] , 
        \q[11][2] , \q[11][1] , \q[11][0] , \q[10][15] , \q[10][14] , 
        \q[10][13] , \q[10][12] , \q[10][11] , \q[10][10] , \q[10][9] , 
        \q[10][8] , \q[10][7] , \q[10][6] , \q[10][5] , \q[10][4] , \q[10][3] , 
        \q[10][2] , \q[10][1] , \q[10][0] , \q[9][15] , \q[9][14] , \q[9][13] , 
        \q[9][12] , \q[9][11] , \q[9][10] , \q[9][9] , \q[9][8] , \q[9][7] , 
        \q[9][6] , \q[9][5] , \q[9][4] , \q[9][3] , \q[9][2] , \q[9][1] , 
        \q[9][0] , \q[8][15] , \q[8][14] , \q[8][13] , \q[8][12] , \q[8][11] , 
        \q[8][10] , \q[8][9] , \q[8][8] , \q[8][7] , \q[8][6] , \q[8][5] , 
        \q[8][4] , \q[8][3] , \q[8][2] , \q[8][1] , \q[8][0] , \q[7][15] , 
        \q[7][14] , \q[7][13] , \q[7][12] , \q[7][11] , \q[7][10] , \q[7][9] , 
        \q[7][8] , \q[7][7] , \q[7][6] , \q[7][5] , \q[7][4] , \q[7][3] , 
        \q[7][2] , \q[7][1] , \q[7][0] , \q[6][15] , \q[6][14] , \q[6][13] , 
        \q[6][12] , \q[6][11] , \q[6][10] , \q[6][9] , \q[6][8] , \q[6][7] , 
        \q[6][6] , \q[6][5] , \q[6][4] , \q[6][3] , \q[6][2] , \q[6][1] , 
        \q[6][0] , \q[5][15] , \q[5][14] , \q[5][13] , \q[5][12] , \q[5][11] , 
        \q[5][10] , \q[5][9] , \q[5][8] , \q[5][7] , \q[5][6] , \q[5][5] , 
        \q[5][4] , \q[5][3] , \q[5][2] , \q[5][1] , \q[5][0] , \q[4][15] , 
        \q[4][14] , \q[4][13] , \q[4][12] , \q[4][11] , \q[4][10] , \q[4][9] , 
        \q[4][8] , \q[4][7] , \q[4][6] , \q[4][5] , \q[4][4] , \q[4][3] , 
        \q[4][2] , \q[4][1] , \q[4][0] , \q[3][15] , \q[3][14] , \q[3][13] , 
        \q[3][12] , \q[3][11] , \q[3][10] , \q[3][9] , \q[3][8] , \q[3][7] , 
        \q[3][6] , \q[3][5] , \q[3][4] , \q[3][3] , \q[3][2] , \q[3][1] , 
        \q[3][0] , \q[2][15] , \q[2][14] , \q[2][13] , \q[2][12] , \q[2][11] , 
        \q[2][10] , \q[2][9] , \q[2][8] , \q[2][7] , \q[2][6] , \q[2][5] , 
        \q[2][4] , \q[2][3] , \q[2][2] , \q[2][1] , \q[2][0] , \q[1][15] , 
        \q[1][14] , \q[1][13] , \q[1][12] , \q[1][11] , \q[1][10] , \q[1][9] , 
        \q[1][8] , \q[1][7] , \q[1][6] , \q[1][5] , \q[1][4] , \q[1][3] , 
        \q[1][2] , \q[1][1] , \q[1][0] , \q[0][15] , \q[0][14] , \q[0][13] , 
        \q[0][12] , \q[0][11] , \q[0][10] , \q[0][9] , \q[0][8] , \q[0][7] , 
        \q[0][6] , \q[0][5] , \q[0][4] , \q[0][3] , \q[0][2] , \q[0][1] , 
        \q[0][0] }), .SEL(rd_addr), .MUX(data_out) );
    MUX21H MX1_0_0 ( .A(\q[0][0] ), .B(data_in[0]), .S(\wren[0] ), .Z(
        \din[0][0] ) );
    MUX21H MX1_0_11 ( .A(\q[11][0] ), .B(data_in[0]), .S(\wren[11] ), .Z(
        \din[11][0] ) );
    MUX21H MX1_8_1 ( .A(\q[1][8] ), .B(data_in[8]), .S(\wren[1] ), .Z(
        \din[1][8] ) );
    MUX21H MX1_15_9 ( .A(\q[9][15] ), .B(data_in[15]), .S(\wren[9] ), .Z(
        \din[9][15] ) );
    MUX21H MX1_12_3 ( .A(\q[3][12] ), .B(data_in[12]), .S(\wren[3] ), .Z(
        \din[3][12] ) );
    MUX21H MX1_14_12 ( .A(\q[12][14] ), .B(data_in[14]), .S(\wren[12] ), .Z(
        \din[12][14] ) );
    MUX21H MX1_5_6 ( .A(\q[6][5] ), .B(data_in[5]), .S(\wren[6] ), .Z(
        \din[6][5] ) );
    MUX21H MX1_6_14 ( .A(\q[14][6] ), .B(data_in[6]), .S(\wren[14] ), .Z(
        \din[14][6] ) );
    MUX21H MX1_1_0 ( .A(\q[0][1] ), .B(data_in[1]), .S(\wren[0] ), .Z(
        \din[0][1] ) );
    MUX21H MX1_4_6 ( .A(\q[6][4] ), .B(data_in[4]), .S(\wren[6] ), .Z(
        \din[6][4] ) );
    MUX21H MX1_1_10 ( .A(\q[10][1] ), .B(data_in[1]), .S(\wren[10] ), .Z(
        \din[10][1] ) );
    MUX21H MX1_0_9 ( .A(\q[9][0] ), .B(data_in[0]), .S(\wren[9] ), .Z(
        \din[9][0] ) );
    MUX21H MX1_4_10 ( .A(\q[10][4] ), .B(data_in[4]), .S(\wren[10] ), .Z(
        \din[10][4] ) );
    MUX21H MX1_14_9 ( .A(\q[9][14] ), .B(data_in[14]), .S(\wren[9] ), .Z(
        \din[9][14] ) );
    MUX21H MX1_7_15 ( .A(\q[15][7] ), .B(data_in[7]), .S(\wren[15] ), .Z(
        \din[15][7] ) );
    MUX21H MX1_15_13 ( .A(\q[13][15] ), .B(data_in[15]), .S(\wren[13] ), .Z(
        \din[13][15] ) );
    MUX21H MX1_9_1 ( .A(\q[1][9] ), .B(data_in[9]), .S(\wren[1] ), .Z(
        \din[1][9] ) );
    MUX21H MX1_8_8 ( .A(\q[8][8] ), .B(data_in[8]), .S(\wren[8] ), .Z(
        \din[8][8] ) );
    MUX21H MX1_13_3 ( .A(\q[3][13] ), .B(data_in[13]), .S(\wren[3] ), .Z(
        \din[3][13] ) );
    MUX21H MX1_15_0 ( .A(\q[0][15] ), .B(data_in[15]), .S(\wren[0] ), .Z(
        \din[0][15] ) );
    MUX21H MX1_10_6 ( .A(\q[6][10] ), .B(data_in[10]), .S(\wren[6] ), .Z(
        \din[6][10] ) );
    MUX21H MX1_1_9 ( .A(\q[9][1] ), .B(data_in[1]), .S(\wren[9] ), .Z(
        \din[9][1] ) );
    MUX21H MX1_2_5 ( .A(\q[5][2] ), .B(data_in[2]), .S(\wren[5] ), .Z(
        \din[5][2] ) );
    MUX21H MX1_8_13 ( .A(\q[13][8] ), .B(data_in[8]), .S(\wren[13] ), .Z(
        \din[13][8] ) );
    MUX21H MX1_2_15 ( .A(\q[15][2] ), .B(data_in[2]), .S(\wren[15] ), .Z(
        \din[15][2] ) );
    MUX21H MX1_7_3 ( .A(\q[3][7] ), .B(data_in[7]), .S(\wren[3] ), .Z(
        \din[3][7] ) );
    MUX21H MX1_10_13 ( .A(\q[13][10] ), .B(data_in[10]), .S(\wren[13] ), .Z(
        \din[13][10] ) );
    MUX21H MX1_5_11 ( .A(\q[11][5] ), .B(data_in[5]), .S(\wren[11] ), .Z(
        \din[11][5] ) );
    MUX21H MX1_6_3 ( .A(\q[3][6] ), .B(data_in[6]), .S(\wren[3] ), .Z(
        \din[3][6] ) );
    MUX21H MX1_3_5 ( .A(\q[5][3] ), .B(data_in[3]), .S(\wren[5] ), .Z(
        \din[5][3] ) );
    MUX21H MX1_3_14 ( .A(\q[14][3] ), .B(data_in[3]), .S(\wren[14] ), .Z(
        \din[14][3] ) );
    MUX21H MX1_9_8 ( .A(\q[8][9] ), .B(data_in[9]), .S(\wren[8] ), .Z(
        \din[8][9] ) );
    MUX21H MX1_9_12 ( .A(\q[12][9] ), .B(data_in[9]), .S(\wren[12] ), .Z(
        \din[12][9] ) );
    MUX21H MX1_11_6 ( .A(\q[6][11] ), .B(data_in[11]), .S(\wren[6] ), .Z(
        \din[6][11] ) );
    MUX21H MX1_14_0 ( .A(\q[0][14] ), .B(data_in[14]), .S(\wren[0] ), .Z(
        \din[0][14] ) );
    MUX21H MX1_9_15 ( .A(\q[15][9] ), .B(data_in[9]), .S(\wren[15] ), .Z(
        \din[15][9] ) );
    MUX21H MX1_11_12 ( .A(\q[12][11] ), .B(data_in[11]), .S(\wren[12] ), .Z(
        \din[12][11] ) );
    MUX21H MX1_14_7 ( .A(\q[7][14] ), .B(data_in[14]), .S(\wren[7] ), .Z(
        \din[7][14] ) );
    MUX21H MX1_11_1 ( .A(\q[1][11] ), .B(data_in[11]), .S(\wren[1] ), .Z(
        \din[1][11] ) );
    MUX21H MX1_3_13 ( .A(\q[13][3] ), .B(data_in[3]), .S(\wren[13] ), .Z(
        \din[13][3] ) );
    MUX21H MX1_11_15 ( .A(\q[15][11] ), .B(data_in[11]), .S(\wren[15] ), .Z(
        \din[15][11] ) );
    MUX21H MX1_4_8 ( .A(\q[8][4] ), .B(data_in[4]), .S(\wren[8] ), .Z(
        \din[8][4] ) );
    MUX21H MX1_3_2 ( .A(\q[2][3] ), .B(data_in[3]), .S(\wren[2] ), .Z(
        \din[2][3] ) );
    MUX21H MX1_6_4 ( .A(\q[4][6] ), .B(data_in[6]), .S(\wren[4] ), .Z(
        \din[4][6] ) );
    MUX21H MX1_2_2 ( .A(\q[2][2] ), .B(data_in[2]), .S(\wren[2] ), .Z(
        \din[2][2] ) );
    MUX21H MX1_2_12 ( .A(\q[12][2] ), .B(data_in[2]), .S(\wren[12] ), .Z(
        \din[12][2] ) );
    MUX21H MX1_5_8 ( .A(\q[8][5] ), .B(data_in[5]), .S(\wren[8] ), .Z(
        \din[8][5] ) );
    MUX21H MX1_8_14 ( .A(\q[14][8] ), .B(data_in[8]), .S(\wren[14] ), .Z(
        \din[14][8] ) );
    MUX21H MX1_10_14 ( .A(\q[14][10] ), .B(data_in[10]), .S(\wren[14] ), .Z(
        \din[14][10] ) );
    MUX21H MX1_7_4 ( .A(\q[4][7] ), .B(data_in[7]), .S(\wren[4] ), .Z(
        \din[4][7] ) );
    MUX21H MX1_7_12 ( .A(\q[12][7] ), .B(data_in[7]), .S(\wren[12] ), .Z(
        \din[12][7] ) );
    MUX21H MX1_10_1 ( .A(\q[1][10] ), .B(data_in[10]), .S(\wren[1] ), .Z(
        \din[1][10] ) );
    MUX21H MX1_15_7 ( .A(\q[7][15] ), .B(data_in[15]), .S(\wren[7] ), .Z(
        \din[7][15] ) );
    MUX21H MX1_9_6 ( .A(\q[6][9] ), .B(data_in[9]), .S(\wren[6] ), .Z(
        \din[6][9] ) );
    MUX21H MX1_11_8 ( .A(\q[8][11] ), .B(data_in[11]), .S(\wren[8] ), .Z(
        \din[8][11] ) );
    MUX21H MX1_13_4 ( .A(\q[4][13] ), .B(data_in[13]), .S(\wren[4] ), .Z(
        \din[4][13] ) );
    MUX21H MX1_15_14 ( .A(\q[14][15] ), .B(data_in[15]), .S(\wren[14] ), .Z(
        \din[14][15] ) );
    MUX21H MX1_0_1 ( .A(\q[1][0] ), .B(data_in[0]), .S(\wren[1] ), .Z(
        \din[1][0] ) );
    MUX21H MX1_0_6 ( .A(\q[6][0] ), .B(data_in[0]), .S(\wren[6] ), .Z(
        \din[6][0] ) );
    MUX21H MX1_0_7 ( .A(\q[7][0] ), .B(data_in[0]), .S(\wren[7] ), .Z(
        \din[7][0] ) );
    MUX21H MX1_1_7 ( .A(\q[7][1] ), .B(data_in[1]), .S(\wren[7] ), .Z(
        \din[7][1] ) );
    MUX21H MX1_4_1 ( .A(\q[1][4] ), .B(data_in[4]), .S(\wren[1] ), .Z(
        \din[1][4] ) );
    MUX21H MX1_13_11 ( .A(\q[11][13] ), .B(data_in[13]), .S(\wren[11] ), .Z(
        \din[11][13] ) );
    MUX21H MX1_5_1 ( .A(\q[1][5] ), .B(data_in[5]), .S(\wren[1] ), .Z(
        \din[1][5] ) );
    MUX21H MX1_6_13 ( .A(\q[13][6] ), .B(data_in[6]), .S(\wren[13] ), .Z(
        \din[13][6] ) );
    MUX21H MX1_14_15 ( .A(\q[15][14] ), .B(data_in[14]), .S(\wren[15] ), .Z(
        \din[15][14] ) );
    MUX21H MX1_8_6 ( .A(\q[6][8] ), .B(data_in[8]), .S(\wren[6] ), .Z(
        \din[6][8] ) );
    MUX21H MX1_8_15 ( .A(\q[15][8] ), .B(data_in[8]), .S(\wren[15] ), .Z(
        \din[15][8] ) );
    MUX21H MX1_10_8 ( .A(\q[8][10] ), .B(data_in[10]), .S(\wren[8] ), .Z(
        \din[8][10] ) );
    MUX21H MX1_12_10 ( .A(\q[10][12] ), .B(data_in[12]), .S(\wren[10] ), .Z(
        \din[10][12] ) );
    MUX21H MX1_12_4 ( .A(\q[4][12] ), .B(data_in[12]), .S(\wren[4] ), .Z(
        \din[4][12] ) );
    MUX21H MX1_10_0 ( .A(\q[0][10] ), .B(data_in[10]), .S(\wren[0] ), .Z(
        \din[0][10] ) );
    MUX21H MX1_15_6 ( .A(\q[6][15] ), .B(data_in[15]), .S(\wren[6] ), .Z(
        \din[6][15] ) );
    MUX21H MX1_2_3 ( .A(\q[3][2] ), .B(data_in[2]), .S(\wren[3] ), .Z(
        \din[3][2] ) );
    MUX21H MX1_2_13 ( .A(\q[13][2] ), .B(data_in[2]), .S(\wren[13] ), .Z(
        \din[13][2] ) );
    MUX21H MX1_5_9 ( .A(\q[9][5] ), .B(data_in[5]), .S(\wren[9] ), .Z(
        \din[9][5] ) );
    MUX21H MX1_7_5 ( .A(\q[5][7] ), .B(data_in[7]), .S(\wren[5] ), .Z(
        \din[5][7] ) );
    MUX21H MX1_10_15 ( .A(\q[15][10] ), .B(data_in[10]), .S(\wren[15] ), .Z(
        \din[15][10] ) );
    MUX21H MX1_4_9 ( .A(\q[9][4] ), .B(data_in[4]), .S(\wren[9] ), .Z(
        \din[9][4] ) );
    MUX21H MX1_3_3 ( .A(\q[3][3] ), .B(data_in[3]), .S(\wren[3] ), .Z(
        \din[3][3] ) );
    MUX21H MX1_6_5 ( .A(\q[5][6] ), .B(data_in[6]), .S(\wren[5] ), .Z(
        \din[5][6] ) );
    MUX21H MX1_9_14 ( .A(\q[14][9] ), .B(data_in[9]), .S(\wren[14] ), .Z(
        \din[14][9] ) );
    MUX21H MX1_14_6 ( .A(\q[6][14] ), .B(data_in[14]), .S(\wren[6] ), .Z(
        \din[6][14] ) );
    MUX21H MX1_11_0 ( .A(\q[0][11] ), .B(data_in[11]), .S(\wren[0] ), .Z(
        \din[0][11] ) );
    MUX21H MX1_3_12 ( .A(\q[12][3] ), .B(data_in[3]), .S(\wren[12] ), .Z(
        \din[12][3] ) );
    MUX21H MX1_11_14 ( .A(\q[14][11] ), .B(data_in[11]), .S(\wren[14] ), .Z(
        \din[14][11] ) );
    MUX21H MX1_5_0 ( .A(\q[0][5] ), .B(data_in[5]), .S(\wren[0] ), .Z(
        \din[0][5] ) );
    MUX21H MX1_8_7 ( .A(\q[7][8] ), .B(data_in[8]), .S(\wren[7] ), .Z(
        \din[7][8] ) );
    MUX21H MX1_10_9 ( .A(\q[9][10] ), .B(data_in[10]), .S(\wren[9] ), .Z(
        \din[9][10] ) );
    MUX21H MX1_12_11 ( .A(\q[11][12] ), .B(data_in[12]), .S(\wren[11] ), .Z(
        \din[11][12] ) );
    MUX21H MX1_12_5 ( .A(\q[5][12] ), .B(data_in[12]), .S(\wren[5] ), .Z(
        \din[5][12] ) );
    MUX21H MX1_6_12 ( .A(\q[12][6] ), .B(data_in[6]), .S(\wren[12] ), .Z(
        \din[12][6] ) );
    MUX21H MX1_14_14 ( .A(\q[14][14] ), .B(data_in[14]), .S(\wren[14] ), .Z(
        \din[14][14] ) );
    MUX21H MX1_1_6 ( .A(\q[6][1] ), .B(data_in[1]), .S(\wren[6] ), .Z(
        \din[6][1] ) );
    MUX21H MX1_4_0 ( .A(\q[0][4] ), .B(data_in[4]), .S(\wren[0] ), .Z(
        \din[0][4] ) );
    MUX21H MX1_7_13 ( .A(\q[13][7] ), .B(data_in[7]), .S(\wren[13] ), .Z(
        \din[13][7] ) );
    MUX21H MX1_13_10 ( .A(\q[10][13] ), .B(data_in[13]), .S(\wren[10] ), .Z(
        \din[10][13] ) );
    MUX21H MX1_11_9 ( .A(\q[9][11] ), .B(data_in[11]), .S(\wren[9] ), .Z(
        \din[9][11] ) );
    MUX21H MX1_9_7 ( .A(\q[7][9] ), .B(data_in[9]), .S(\wren[7] ), .Z(
        \din[7][9] ) );
    MUX21H MX1_13_5 ( .A(\q[5][13] ), .B(data_in[13]), .S(\wren[5] ), .Z(
        \din[5][13] ) );
    MUX21H MX1_15_15 ( .A(\q[15][15] ), .B(data_in[15]), .S(\wren[15] ), .Z(
        \din[15][15] ) );
    MUX21H MX1_7_14 ( .A(\q[14][7] ), .B(data_in[7]), .S(\wren[14] ), .Z(
        \din[14][7] ) );
    MUX21H MX1_9_0 ( .A(\q[0][9] ), .B(data_in[9]), .S(\wren[0] ), .Z(
        \din[0][9] ) );
    MUX21H MX1_14_8 ( .A(\q[8][14] ), .B(data_in[14]), .S(\wren[8] ), .Z(
        \din[8][14] ) );
    MUX21H MX1_15_12 ( .A(\q[12][15] ), .B(data_in[15]), .S(\wren[12] ), .Z(
        \din[12][15] ) );
    MUX21H MX1_13_2 ( .A(\q[2][13] ), .B(data_in[13]), .S(\wren[2] ), .Z(
        \din[2][13] ) );
    MUX21H MX1_1_1 ( .A(\q[1][1] ), .B(data_in[1]), .S(\wren[1] ), .Z(
        \din[1][1] ) );
    MUX21H MX1_1_11 ( .A(\q[11][1] ), .B(data_in[1]), .S(\wren[11] ), .Z(
        \din[11][1] ) );
    MUX21H MX1_4_7 ( .A(\q[7][4] ), .B(data_in[4]), .S(\wren[7] ), .Z(
        \din[7][4] ) );
    MUX21H MX1_14_13 ( .A(\q[13][14] ), .B(data_in[14]), .S(\wren[13] ), .Z(
        \din[13][14] ) );
    MUX21H MX1_0_2 ( .A(\q[2][0] ), .B(data_in[0]), .S(\wren[2] ), .Z(
        \din[2][0] ) );
    MUX21H MX1_0_3 ( .A(\q[3][0] ), .B(data_in[0]), .S(\wren[3] ), .Z(
        \din[3][0] ) );
    MUX21H MX1_0_8 ( .A(\q[8][0] ), .B(data_in[0]), .S(\wren[8] ), .Z(
        \din[8][0] ) );
    MUX21H MX1_0_10 ( .A(\q[10][0] ), .B(data_in[0]), .S(\wren[10] ), .Z(
        \din[10][0] ) );
    MUX21H MX1_5_7 ( .A(\q[7][5] ), .B(data_in[5]), .S(\wren[7] ), .Z(
        \din[7][5] ) );
    MUX21H MX1_6_15 ( .A(\q[15][6] ), .B(data_in[6]), .S(\wren[15] ), .Z(
        \din[15][6] ) );
    MUX21H MX1_8_0 ( .A(\q[0][8] ), .B(data_in[8]), .S(\wren[0] ), .Z(
        \din[0][8] ) );
    MUX21H MX1_1_8 ( .A(\q[8][1] ), .B(data_in[1]), .S(\wren[8] ), .Z(
        \din[8][1] ) );
    MUX21H MX1_3_15 ( .A(\q[15][3] ), .B(data_in[3]), .S(\wren[15] ), .Z(
        \din[15][3] ) );
    MUX21H MX1_12_2 ( .A(\q[2][12] ), .B(data_in[12]), .S(\wren[2] ), .Z(
        \din[2][12] ) );
    MUX21H MX1_15_8 ( .A(\q[8][15] ), .B(data_in[15]), .S(\wren[8] ), .Z(
        \din[8][15] ) );
    MUX21H MX1_9_9 ( .A(\q[9][9] ), .B(data_in[9]), .S(\wren[9] ), .Z(
        \din[9][9] ) );
    MUX21H MX1_11_7 ( .A(\q[7][11] ), .B(data_in[11]), .S(\wren[7] ), .Z(
        \din[7][11] ) );
    MUX21H MX1_9_13 ( .A(\q[13][9] ), .B(data_in[9]), .S(\wren[13] ), .Z(
        \din[13][9] ) );
    MUX21H MX1_14_1 ( .A(\q[1][14] ), .B(data_in[14]), .S(\wren[1] ), .Z(
        \din[1][14] ) );
    MUX21H MX1_11_13 ( .A(\q[13][11] ), .B(data_in[11]), .S(\wren[13] ), .Z(
        \din[13][11] ) );
    MUX21H MX1_5_10 ( .A(\q[10][5] ), .B(data_in[5]), .S(\wren[10] ), .Z(
        \din[10][5] ) );
    MUX21H MX1_6_2 ( .A(\q[2][6] ), .B(data_in[6]), .S(\wren[2] ), .Z(
        \din[2][6] ) );
    MUX21H MX1_3_4 ( .A(\q[4][3] ), .B(data_in[3]), .S(\wren[4] ), .Z(
        \din[4][3] ) );
    MUX21H MX1_0_12 ( .A(\q[12][0] ), .B(data_in[0]), .S(\wren[12] ), .Z(
        \din[12][0] ) );
    MUX21H MX1_2_4 ( .A(\q[4][2] ), .B(data_in[2]), .S(\wren[4] ), .Z(
        \din[4][2] ) );
    MUX21H MX1_8_12 ( .A(\q[12][8] ), .B(data_in[8]), .S(\wren[12] ), .Z(
        \din[12][8] ) );
    MUX21H MX1_2_14 ( .A(\q[14][2] ), .B(data_in[2]), .S(\wren[14] ), .Z(
        \din[14][2] ) );
    MUX21H MX1_7_2 ( .A(\q[2][7] ), .B(data_in[7]), .S(\wren[2] ), .Z(
        \din[2][7] ) );
    MUX21H MX1_4_11 ( .A(\q[11][4] ), .B(data_in[4]), .S(\wren[11] ), .Z(
        \din[11][4] ) );
    MUX21H MX1_10_12 ( .A(\q[12][10] ), .B(data_in[10]), .S(\wren[12] ), .Z(
        \din[12][10] ) );
    MUX21H MX1_8_9 ( .A(\q[9][8] ), .B(data_in[8]), .S(\wren[9] ), .Z(
        \din[9][8] ) );
    MUX21H MX1_10_7 ( .A(\q[7][10] ), .B(data_in[10]), .S(\wren[7] ), .Z(
        \din[7][10] ) );
    MUX21H MX1_15_1 ( .A(\q[1][15] ), .B(data_in[15]), .S(\wren[1] ), .Z(
        \din[1][15] ) );
    MUX21H MX1_12_0 ( .A(\q[0][12] ), .B(data_in[12]), .S(\wren[0] ), .Z(
        \din[0][12] ) );
    MUX21H MX1_8_2 ( .A(\q[2][8] ), .B(data_in[8]), .S(\wren[2] ), .Z(
        \din[2][8] ) );
    MUX21H MX1_12_14 ( .A(\q[14][12] ), .B(data_in[12]), .S(\wren[14] ), .Z(
        \din[14][12] ) );
    MUX21H MX1_7_9 ( .A(\q[9][7] ), .B(data_in[7]), .S(\wren[9] ), .Z(
        \din[9][7] ) );
    MUX21H MX1_5_5 ( .A(\q[5][5] ), .B(data_in[5]), .S(\wren[5] ), .Z(
        \din[5][5] ) );
    MUX21H MX1_1_3 ( .A(\q[3][1] ), .B(data_in[1]), .S(\wren[3] ), .Z(
        \din[3][1] ) );
    MUX21H MX1_6_9 ( .A(\q[9][6] ), .B(data_in[6]), .S(\wren[9] ), .Z(
        \din[9][6] ) );
    MUX21H MX1_14_11 ( .A(\q[11][14] ), .B(data_in[14]), .S(\wren[11] ), .Z(
        \din[11][14] ) );
    MUX21H MX1_1_13 ( .A(\q[13][1] ), .B(data_in[1]), .S(\wren[13] ), .Z(
        \din[13][1] ) );
    MUX21H MX1_2_1 ( .A(\q[1][2] ), .B(data_in[2]), .S(\wren[1] ), .Z(
        \din[1][2] ) );
    MUX21H MX1_2_6 ( .A(\q[6][2] ), .B(data_in[2]), .S(\wren[6] ), .Z(
        \din[6][2] ) );
    MUX21H MX1_4_5 ( .A(\q[5][4] ), .B(data_in[4]), .S(\wren[5] ), .Z(
        \din[5][4] ) );
    MUX21H MX1_13_15 ( .A(\q[15][13] ), .B(data_in[13]), .S(\wren[15] ), .Z(
        \din[15][13] ) );
    MUX21H MX1_4_13 ( .A(\q[13][4] ), .B(data_in[4]), .S(\wren[13] ), .Z(
        \din[13][4] ) );
    MUX21H MX1_9_2 ( .A(\q[2][9] ), .B(data_in[9]), .S(\wren[2] ), .Z(
        \din[2][9] ) );
    MUX21H MX1_13_0 ( .A(\q[0][13] ), .B(data_in[13]), .S(\wren[0] ), .Z(
        \din[0][13] ) );
    MUX21H MX1_15_10 ( .A(\q[10][15] ), .B(data_in[15]), .S(\wren[10] ), .Z(
        \din[10][15] ) );
    MUX21H MX1_12_9 ( .A(\q[9][12] ), .B(data_in[12]), .S(\wren[9] ), .Z(
        \din[9][12] ) );
    MUX21H MX1_7_0 ( .A(\q[0][7] ), .B(data_in[7]), .S(\wren[0] ), .Z(
        \din[0][7] ) );
    MUX21H MX1_10_5 ( .A(\q[5][10] ), .B(data_in[10]), .S(\wren[5] ), .Z(
        \din[5][10] ) );
    MUX21H MX1_15_3 ( .A(\q[3][15] ), .B(data_in[15]), .S(\wren[3] ), .Z(
        \din[3][15] ) );
    MUX21H MX1_10_10 ( .A(\q[10][10] ), .B(data_in[10]), .S(\wren[10] ), .Z(
        \din[10][10] ) );
    MUX21H MX1_8_10 ( .A(\q[10][8] ), .B(data_in[8]), .S(\wren[10] ), .Z(
        \din[10][8] ) );
    MUX21H MX1_3_6 ( .A(\q[6][3] ), .B(data_in[3]), .S(\wren[6] ), .Z(
        \din[6][3] ) );
    MUX21H MX1_3_10 ( .A(\q[10][3] ), .B(data_in[3]), .S(\wren[10] ), .Z(
        \din[10][3] ) );
    MUX21H MX1_5_12 ( .A(\q[12][5] ), .B(data_in[5]), .S(\wren[12] ), .Z(
        \din[12][5] ) );
    MUX21H MX1_6_0 ( .A(\q[0][6] ), .B(data_in[6]), .S(\wren[0] ), .Z(
        \din[0][6] ) );
    MUX21H MX1_9_11 ( .A(\q[11][9] ), .B(data_in[9]), .S(\wren[11] ), .Z(
        \din[11][9] ) );
    MUX21H MX1_11_11 ( .A(\q[11][11] ), .B(data_in[11]), .S(\wren[11] ), .Z(
        \din[11][11] ) );
    MUX21H MX1_13_9 ( .A(\q[9][13] ), .B(data_in[13]), .S(\wren[9] ), .Z(
        \din[9][13] ) );
    MUX21H MX1_14_3 ( .A(\q[3][14] ), .B(data_in[14]), .S(\wren[3] ), .Z(
        \din[3][14] ) );
    MUX21H MX1_11_5 ( .A(\q[5][11] ), .B(data_in[11]), .S(\wren[5] ), .Z(
        \din[5][11] ) );
    MUX21H MX1_3_1 ( .A(\q[1][3] ), .B(data_in[3]), .S(\wren[1] ), .Z(
        \din[1][3] ) );
    MUX21H MX1_5_15 ( .A(\q[15][5] ), .B(data_in[5]), .S(\wren[15] ), .Z(
        \din[15][5] ) );
    MUX21H MX1_6_7 ( .A(\q[7][6] ), .B(data_in[6]), .S(\wren[7] ), .Z(
        \din[7][6] ) );
    MUX21H MX1_11_2 ( .A(\q[2][11] ), .B(data_in[11]), .S(\wren[2] ), .Z(
        \din[2][11] ) );
    MUX21H MX1_14_4 ( .A(\q[4][14] ), .B(data_in[14]), .S(\wren[4] ), .Z(
        \din[4][14] ) );
    MUX21H MX1_2_11 ( .A(\q[11][2] ), .B(data_in[2]), .S(\wren[11] ), .Z(
        \din[11][2] ) );
    MUX21H MX1_3_8 ( .A(\q[8][3] ), .B(data_in[3]), .S(\wren[8] ), .Z(
        \din[8][3] ) );
    MUX21H MX1_4_14 ( .A(\q[14][4] ), .B(data_in[4]), .S(\wren[14] ), .Z(
        \din[14][4] ) );
    MUX21H MX1_7_7 ( .A(\q[7][7] ), .B(data_in[7]), .S(\wren[7] ), .Z(
        \din[7][7] ) );
    MUX21H MX1_10_2 ( .A(\q[2][10] ), .B(data_in[10]), .S(\wren[2] ), .Z(
        \din[2][10] ) );
    MUX21H MX1_15_4 ( .A(\q[4][15] ), .B(data_in[15]), .S(\wren[4] ), .Z(
        \din[4][15] ) );
    MUX21H MX1_13_7 ( .A(\q[7][13] ), .B(data_in[13]), .S(\wren[7] ), .Z(
        \din[7][13] ) );
    MUX21H MX1_7_11 ( .A(\q[11][7] ), .B(data_in[7]), .S(\wren[11] ), .Z(
        \din[11][7] ) );
    MUX21H MX1_9_5 ( .A(\q[5][9] ), .B(data_in[9]), .S(\wren[5] ), .Z(
        \din[5][9] ) );
    MUX21H MX1_4_2 ( .A(\q[2][4] ), .B(data_in[4]), .S(\wren[2] ), .Z(
        \din[2][4] ) );
    MUX21H MX1_13_12 ( .A(\q[12][13] ), .B(data_in[13]), .S(\wren[12] ), .Z(
        \din[12][13] ) );
    MUX21H MX1_0_4 ( .A(\q[4][0] ), .B(data_in[0]), .S(\wren[4] ), .Z(
        \din[4][0] ) );
    MUX21H MX1_1_4 ( .A(\q[4][1] ), .B(data_in[1]), .S(\wren[4] ), .Z(
        \din[4][1] ) );
    MUX21H MX1_1_14 ( .A(\q[14][1] ), .B(data_in[1]), .S(\wren[14] ), .Z(
        \din[14][1] ) );
    MUX21H MX1_2_8 ( .A(\q[8][2] ), .B(data_in[2]), .S(\wren[8] ), .Z(
        \din[8][2] ) );
    MUX21H MX1_0_5 ( .A(\q[5][0] ), .B(data_in[0]), .S(\wren[5] ), .Z(
        \din[5][0] ) );
    MUX21H MX1_0_14 ( .A(\q[14][0] ), .B(data_in[0]), .S(\wren[14] ), .Z(
        \din[14][0] ) );
    MUX21H MX1_0_15 ( .A(\q[15][0] ), .B(data_in[0]), .S(\wren[15] ), .Z(
        \din[15][0] ) );
    MUX21H MX1_5_2 ( .A(\q[2][5] ), .B(data_in[5]), .S(\wren[2] ), .Z(
        \din[2][5] ) );
    MUX21H MX1_6_10 ( .A(\q[10][6] ), .B(data_in[6]), .S(\wren[10] ), .Z(
        \din[10][6] ) );
    MUX21H MX1_8_5 ( .A(\q[5][8] ), .B(data_in[8]), .S(\wren[5] ), .Z(
        \din[5][8] ) );
    MUX21H MX1_12_7 ( .A(\q[7][12] ), .B(data_in[12]), .S(\wren[7] ), .Z(
        \din[7][12] ) );
    MUX21H MX1_12_13 ( .A(\q[13][12] ), .B(data_in[12]), .S(\wren[13] ), .Z(
        \din[13][12] ) );
    MUX21H MX1_2_0 ( .A(\q[0][2] ), .B(data_in[2]), .S(\wren[0] ), .Z(
        \din[0][2] ) );
    MUX21H MX1_2_10 ( .A(\q[10][2] ), .B(data_in[2]), .S(\wren[10] ), .Z(
        \din[10][2] ) );
    MUX21H MX1_4_15 ( .A(\q[15][4] ), .B(data_in[4]), .S(\wren[15] ), .Z(
        \din[15][4] ) );
    MUX21H MX1_10_3 ( .A(\q[3][10] ), .B(data_in[10]), .S(\wren[3] ), .Z(
        \din[3][10] ) );
    MUX21H MX1_15_5 ( .A(\q[5][15] ), .B(data_in[15]), .S(\wren[5] ), .Z(
        \din[5][15] ) );
    MUX21H MX1_3_0 ( .A(\q[0][3] ), .B(data_in[3]), .S(\wren[0] ), .Z(
        \din[0][3] ) );
    MUX21H MX1_5_14 ( .A(\q[14][5] ), .B(data_in[5]), .S(\wren[14] ), .Z(
        \din[14][5] ) );
    MUX21H MX1_6_6 ( .A(\q[6][6] ), .B(data_in[6]), .S(\wren[6] ), .Z(
        \din[6][6] ) );
    MUX21H MX1_7_6 ( .A(\q[6][7] ), .B(data_in[7]), .S(\wren[6] ), .Z(
        \din[6][7] ) );
    MUX21H MX1_3_11 ( .A(\q[11][3] ), .B(data_in[3]), .S(\wren[11] ), .Z(
        \din[11][3] ) );
    MUX21H MX1_11_3 ( .A(\q[3][11] ), .B(data_in[11]), .S(\wren[3] ), .Z(
        \din[3][11] ) );
    MUX21H MX1_12_6 ( .A(\q[6][12] ), .B(data_in[12]), .S(\wren[6] ), .Z(
        \din[6][12] ) );
    MUX21H MX1_14_5 ( .A(\q[5][14] ), .B(data_in[14]), .S(\wren[5] ), .Z(
        \din[5][14] ) );
    MUX21H MX1_8_4 ( .A(\q[4][8] ), .B(data_in[8]), .S(\wren[4] ), .Z(
        \din[4][8] ) );
    MUX21H MX1_12_12 ( .A(\q[12][12] ), .B(data_in[12]), .S(\wren[12] ), .Z(
        \din[12][12] ) );
    MUX21H MX1_2_9 ( .A(\q[9][2] ), .B(data_in[2]), .S(\wren[9] ), .Z(
        \din[9][2] ) );
    MUX21H MX1_3_9 ( .A(\q[9][3] ), .B(data_in[3]), .S(\wren[9] ), .Z(
        \din[9][3] ) );
    MUX21H MX1_5_3 ( .A(\q[3][5] ), .B(data_in[5]), .S(\wren[3] ), .Z(
        \din[3][5] ) );
    MUX21H MX1_6_11 ( .A(\q[11][6] ), .B(data_in[6]), .S(\wren[11] ), .Z(
        \din[11][6] ) );
    MUX21H MX1_4_3 ( .A(\q[3][4] ), .B(data_in[4]), .S(\wren[3] ), .Z(
        \din[3][4] ) );
    MUX21H MX1_13_13 ( .A(\q[13][13] ), .B(data_in[13]), .S(\wren[13] ), .Z(
        \din[13][13] ) );
    MUX21H MX1_1_2 ( .A(\q[2][1] ), .B(data_in[1]), .S(\wren[2] ), .Z(
        \din[2][1] ) );
    MUX21H MX1_1_5 ( .A(\q[5][1] ), .B(data_in[1]), .S(\wren[5] ), .Z(
        \din[5][1] ) );
    MUX21H MX1_1_12 ( .A(\q[12][1] ), .B(data_in[1]), .S(\wren[12] ), .Z(
        \din[12][1] ) );
    MUX21H MX1_1_15 ( .A(\q[15][1] ), .B(data_in[1]), .S(\wren[15] ), .Z(
        \din[15][1] ) );
    MUX21H MX1_6_8 ( .A(\q[8][6] ), .B(data_in[6]), .S(\wren[8] ), .Z(
        \din[8][6] ) );
    MUX21H MX1_13_6 ( .A(\q[6][13] ), .B(data_in[13]), .S(\wren[6] ), .Z(
        \din[6][13] ) );
    MUX21H MX1_7_10 ( .A(\q[10][7] ), .B(data_in[7]), .S(\wren[10] ), .Z(
        \din[10][7] ) );
    MUX21H MX1_9_3 ( .A(\q[3][9] ), .B(data_in[9]), .S(\wren[3] ), .Z(
        \din[3][9] ) );
    MUX21H MX1_9_4 ( .A(\q[4][9] ), .B(data_in[9]), .S(\wren[4] ), .Z(
        \din[4][9] ) );
    MUX21H MX1_13_1 ( .A(\q[1][13] ), .B(data_in[13]), .S(\wren[1] ), .Z(
        \din[1][13] ) );
    MUX21H MX1_15_11 ( .A(\q[11][15] ), .B(data_in[15]), .S(\wren[11] ), .Z(
        \din[11][15] ) );
    MUX21H MX1_4_4 ( .A(\q[4][4] ), .B(data_in[4]), .S(\wren[4] ), .Z(
        \din[4][4] ) );
    MUX21H MX1_13_14 ( .A(\q[14][13] ), .B(data_in[13]), .S(\wren[14] ), .Z(
        \din[14][13] ) );
    MUX21H MX1_7_8 ( .A(\q[8][7] ), .B(data_in[7]), .S(\wren[8] ), .Z(
        \din[8][7] ) );
    MUX21H MX1_5_4 ( .A(\q[4][5] ), .B(data_in[5]), .S(\wren[4] ), .Z(
        \din[4][5] ) );
    MUX21H MX1_14_10 ( .A(\q[10][14] ), .B(data_in[14]), .S(\wren[10] ), .Z(
        \din[10][14] ) );
    MUX21H MX1_0_13 ( .A(\q[13][0] ), .B(data_in[0]), .S(\wren[13] ), .Z(
        \din[13][0] ) );
    MUX21H MX1_12_1 ( .A(\q[1][12] ), .B(data_in[12]), .S(\wren[1] ), .Z(
        \din[1][12] ) );
    MUX21H MX1_8_3 ( .A(\q[3][8] ), .B(data_in[8]), .S(\wren[3] ), .Z(
        \din[3][8] ) );
    MUX21H MX1_9_10 ( .A(\q[10][9] ), .B(data_in[9]), .S(\wren[10] ), .Z(
        \din[10][9] ) );
    MUX21H MX1_11_10 ( .A(\q[10][11] ), .B(data_in[11]), .S(\wren[10] ), .Z(
        \din[10][11] ) );
    MUX21H MX1_12_15 ( .A(\q[15][12] ), .B(data_in[12]), .S(\wren[15] ), .Z(
        \din[15][12] ) );
    MUX21H MX1_13_8 ( .A(\q[8][13] ), .B(data_in[13]), .S(\wren[8] ), .Z(
        \din[8][13] ) );
    MUX21H MX1_14_2 ( .A(\q[2][14] ), .B(data_in[14]), .S(\wren[2] ), .Z(
        \din[2][14] ) );
    MUX21H MX1_11_4 ( .A(\q[4][11] ), .B(data_in[11]), .S(\wren[4] ), .Z(
        \din[4][11] ) );
    MUX21H MX1_2_7 ( .A(\q[7][2] ), .B(data_in[2]), .S(\wren[7] ), .Z(
        \din[7][2] ) );
    MUX21H MX1_3_7 ( .A(\q[7][3] ), .B(data_in[3]), .S(\wren[7] ), .Z(
        \din[7][3] ) );
    MUX21H MX1_5_13 ( .A(\q[13][5] ), .B(data_in[5]), .S(\wren[13] ), .Z(
        \din[13][5] ) );
    MUX21H MX1_6_1 ( .A(\q[1][6] ), .B(data_in[6]), .S(\wren[1] ), .Z(
        \din[1][6] ) );
    MUX21H MX1_7_1 ( .A(\q[1][7] ), .B(data_in[7]), .S(\wren[1] ), .Z(
        \din[1][7] ) );
    MUX21H MX1_10_11 ( .A(\q[11][10] ), .B(data_in[10]), .S(\wren[11] ), .Z(
        \din[11][10] ) );
    MUX21H MX1_4_12 ( .A(\q[12][4] ), .B(data_in[4]), .S(\wren[12] ), .Z(
        \din[12][4] ) );
    MUX21H MX1_8_11 ( .A(\q[11][8] ), .B(data_in[8]), .S(\wren[11] ), .Z(
        \din[11][8] ) );
    MUX21H MX1_12_8 ( .A(\q[8][12] ), .B(data_in[12]), .S(\wren[8] ), .Z(
        \din[8][12] ) );
    MUX21H MX1_10_4 ( .A(\q[4][10] ), .B(data_in[10]), .S(\wren[4] ), .Z(
        \din[4][10] ) );
    MUX21H MX1_15_2 ( .A(\q[2][15] ), .B(data_in[15]), .S(\wren[2] ), .Z(
        \din[2][15] ) );
    LD1 F0_11_13 ( .D(\din[13][11] ), .G(n73), .Q(\q[13][11] ) );
    LD1 F0_14_2 ( .D(\din[2][14] ), .G(n73), .Q(\q[2][14] ) );
    LD1 F0_9_10 ( .D(\din[10][9] ), .G(n73), .Q(\q[10][9] ) );
    LD1 F0_11_4 ( .D(\din[4][11] ), .G(n73), .Q(\q[4][11] ) );
    LD1 F0_5_13 ( .D(\din[13][5] ), .G(n73), .Q(\q[13][5] ) );
    LD1 F0_3_0 ( .D(\din[0][3] ), .G(n73), .Q(\q[0][3] ) );
    LD1 F0_13_8 ( .D(\din[8][13] ), .G(n73), .Q(\q[8][13] ) );
    LD1 F0_15_2 ( .D(\din[2][15] ), .G(n73), .Q(\q[2][15] ) );
    LD1 F0_10_4 ( .D(\din[4][10] ), .G(n73), .Q(\q[4][10] ) );
    LD1 F0_6_6 ( .D(\din[6][6] ), .G(n73), .Q(\q[6][6] ) );
    LD1 F0_10_12 ( .D(\din[12][10] ), .G(n73), .Q(\q[12][10] ) );
    LD1 F0_7_6 ( .D(\din[6][7] ), .G(n73), .Q(\q[6][7] ) );
    LD1 F0_12_8 ( .D(\din[8][12] ), .G(n73), .Q(\q[8][12] ) );
    LD1 F0_8_11 ( .D(\din[11][8] ), .G(n73), .Q(\q[11][8] ) );
    LD1 F0_4_12 ( .D(\din[12][4] ), .G(n73), .Q(\q[12][4] ) );
    LD1 F0_2_0 ( .D(\din[0][2] ), .G(n73), .Q(\q[0][2] ) );
    LD1 F0_9_4 ( .D(\din[4][9] ), .G(n73), .Q(\q[4][9] ) );
    LD1 F0_1_12 ( .D(\din[12][1] ), .G(n73), .Q(\q[12][1] ) );
    LD1 F0_15_12 ( .D(\din[12][15] ), .G(n73), .Q(\q[12][15] ) );
    LD1 F0_13_1 ( .D(\din[1][13] ), .G(n73), .Q(\q[1][13] ) );
    LD1 F0_4_3 ( .D(\din[3][4] ), .G(n73), .Q(\q[3][4] ) );
    LD1 F0_5_3 ( .D(\din[3][5] ), .G(n73), .Q(\q[3][5] ) );
    LD1 F0_3_9 ( .D(\din[9][3] ), .G(n73), .Q(\q[9][3] ) );
    LD1 F0_1_5 ( .D(\din[5][1] ), .G(n73), .Q(\q[5][1] ) );
    LD1 F0_0_13 ( .D(\din[13][0] ), .G(n73), .Q(\q[13][0] ) );
    LD1 F0_14_13 ( .D(\din[13][14] ), .G(n73), .Q(\q[13][14] ) );
    LD1 F0_12_1 ( .D(\din[1][12] ), .G(n73), .Q(\q[1][12] ) );
    LD1 F0_8_4 ( .D(\din[4][8] ), .G(n73), .Q(\q[4][8] ) );
    LD1 F0_12_11 ( .D(\din[11][12] ), .G(n73), .Q(\q[11][12] ) );
    LD1 F0_8_3 ( .D(\din[3][8] ), .G(n73), .Q(\q[3][8] ) );
    LD1 F0_6_11 ( .D(\din[11][6] ), .G(n73), .Q(\q[11][6] ) );
    LD1 F0_2_9 ( .D(\din[9][2] ), .G(n73), .Q(\q[9][2] ) );
    LD1 F0_14_14 ( .D(\din[14][14] ), .G(n73), .Q(\q[14][14] ) );
    LD1 F0_0_5 ( .D(\din[5][0] ), .G(n73), .Q(\q[5][0] ) );
    LD1 F0_7_8 ( .D(\din[8][7] ), .G(n73), .Q(\q[8][7] ) );
    LD1 F0_5_4 ( .D(\din[4][5] ), .G(n73), .Q(\q[4][5] ) );
    LD1 F0_13_10 ( .D(\din[10][13] ), .G(n73), .Q(\q[10][13] ) );
    LD1 F0_12_6 ( .D(\din[6][12] ), .G(n73), .Q(\q[6][12] ) );
    LD1 F0_4_4 ( .D(\din[4][4] ), .G(n73), .Q(\q[4][4] ) );
    LD1 F0_7_10 ( .D(\din[10][7] ), .G(n73), .Q(\q[10][7] ) );
    LD1 F0_1_2 ( .D(\din[2][1] ), .G(n73), .Q(\q[2][1] ) );
    LD1 F0_0_14 ( .D(\din[14][0] ), .G(n73), .Q(\q[14][0] ) );
    LD1 F0_13_6 ( .D(\din[6][13] ), .G(n73), .Q(\q[6][13] ) );
    LD1 F0_15_15 ( .D(\din[15][15] ), .G(n73), .Q(\q[15][15] ) );
    LD1 F0_6_8 ( .D(\din[8][6] ), .G(n73), .Q(\q[8][6] ) );
    LD1 F0_9_3 ( .D(\din[3][9] ), .G(n73), .Q(\q[3][9] ) );
    LD1 F0_15_5 ( .D(\din[5][15] ), .G(n73), .Q(\q[5][15] ) );
    LD1 F0_10_3 ( .D(\din[3][10] ), .G(n73), .Q(\q[3][10] ) );
    LD1 F0_4_15 ( .D(\din[15][4] ), .G(n73), .Q(\q[15][4] ) );
    LD1 F0_2_10 ( .D(\din[10][2] ), .G(n73), .Q(\q[10][2] ) );
    LD1 F0_10_15 ( .D(\din[15][10] ), .G(n73), .Q(\q[15][10] ) );
    LD1 F0_7_1 ( .D(\din[1][7] ), .G(n73), .Q(\q[1][7] ) );
    LD1 F0_14_5 ( .D(\din[5][14] ), .G(n73), .Q(\q[5][14] ) );
    LD1 F0_11_3 ( .D(\din[3][11] ), .G(n73), .Q(\q[3][11] ) );
    LD1 F0_6_1 ( .D(\din[1][6] ), .G(n73), .Q(\q[1][6] ) );
    LD1 F0_3_11 ( .D(\din[11][3] ), .G(n73), .Q(\q[11][3] ) );
    LD1 F0_2_7 ( .D(\din[7][2] ), .G(n73), .Q(\q[7][2] ) );
    LD1 F0_11_14 ( .D(\din[14][11] ), .G(n73), .Q(\q[14][11] ) );
    LD1 F0_5_14 ( .D(\din[14][5] ), .G(n73), .Q(\q[14][5] ) );
    LD1 F0_15_14 ( .D(\din[14][15] ), .G(n73), .Q(\q[14][15] ) );
    LD1 F0_3_7 ( .D(\din[7][3] ), .G(n73), .Q(\q[7][3] ) );
    LD1 F0_1_15 ( .D(\din[15][1] ), .G(n73), .Q(\q[15][1] ) );
    LD1 F0_9_2 ( .D(\din[2][9] ), .G(n73), .Q(\q[2][9] ) );
    LD1 F0_13_11 ( .D(\din[11][13] ), .G(n73), .Q(\q[11][13] ) );
    LD1 F0_4_5 ( .D(\din[5][4] ), .G(n73), .Q(\q[5][4] ) );
    LD1 F0_1_14 ( .D(\din[14][1] ), .G(n73), .Q(\q[14][1] ) );
    LD1 F0_1_3 ( .D(\din[3][1] ), .G(n73), .Q(\q[3][1] ) );
    LD1 F0_13_7 ( .D(\din[7][13] ), .G(n73), .Q(\q[7][13] ) );
    LD1 F0_7_11 ( .D(\din[11][7] ), .G(n73), .Q(\q[11][7] ) );
    LD1 F0_6_9 ( .D(\din[9][6] ), .G(n73), .Q(\q[9][6] ) );
    LD1 F0_14_15 ( .D(\din[15][14] ), .G(n73), .Q(\q[15][14] ) );
    LD1 F0_12_7 ( .D(\din[7][12] ), .G(n73), .Q(\q[7][12] ) );
    LD1 F0_7_9 ( .D(\din[9][7] ), .G(n73), .Q(\q[9][7] ) );
    LD1 F0_5_5 ( .D(\din[5][5] ), .G(n73), .Q(\q[5][5] ) );
    LD1 F0_12_10 ( .D(\din[10][12] ), .G(n73), .Q(\q[10][12] ) );
    LD1 F0_8_2 ( .D(\din[2][8] ), .G(n73), .Q(\q[2][8] ) );
    LD1 F0_6_10 ( .D(\din[10][6] ), .G(n73), .Q(\q[10][6] ) );
    LD1 F0_11_15 ( .D(\din[15][11] ), .G(n73), .Q(\q[15][11] ) );
    LD1 F0_5_15 ( .D(\din[15][5] ), .G(n73), .Q(\q[15][5] ) );
    LD1 F0_14_4 ( .D(\din[4][14] ), .G(n73), .Q(\q[4][14] ) );
    LD1 F0_11_2 ( .D(\din[2][11] ), .G(n73), .Q(\q[2][11] ) );
    LD1 F0_6_0 ( .D(\din[0][6] ), .G(n73), .Q(\q[0][6] ) );
    LD1 F0_3_10 ( .D(\din[10][3] ), .G(n73), .Q(\q[10][3] ) );
    LD1 F0_3_6 ( .D(\din[6][3] ), .G(n73), .Q(\q[6][3] ) );
    LD1 F0_15_4 ( .D(\din[4][15] ), .G(n73), .Q(\q[4][15] ) );
    LD1 F0_10_2 ( .D(\din[2][10] ), .G(n73), .Q(\q[2][10] ) );
    LD1 F0_4_14 ( .D(\din[14][4] ), .G(n73), .Q(\q[14][4] ) );
    LD1 F0_7_0 ( .D(\din[0][7] ), .G(n73), .Q(\q[0][7] ) );
    LD1 F0_10_14 ( .D(\din[14][10] ), .G(n73), .Q(\q[14][10] ) );
    LD1 F0_15_3 ( .D(\din[3][15] ), .G(n73), .Q(\q[3][15] ) );
    LD1 F0_10_13 ( .D(\din[13][10] ), .G(n73), .Q(\q[13][10] ) );
    LD1 F0_10_5 ( .D(\din[5][10] ), .G(n73), .Q(\q[5][10] ) );
    LD1 F0_8_10 ( .D(\din[10][8] ), .G(n73), .Q(\q[10][8] ) );
    LD1 F0_12_9 ( .D(\din[9][12] ), .G(n73), .Q(\q[9][12] ) );
    LD1 F0_7_7 ( .D(\din[7][7] ), .G(n73), .Q(\q[7][7] ) );
    LD1 F0_2_11 ( .D(\din[11][2] ), .G(n73), .Q(\q[11][2] ) );
    LD1 F0_2_6 ( .D(\din[6][2] ), .G(n73), .Q(\q[6][2] ) );
    LD1 F0_14_3 ( .D(\din[3][14] ), .G(n73), .Q(\q[3][14] ) );
    LD1 F0_9_11 ( .D(\din[11][9] ), .G(n73), .Q(\q[11][9] ) );
    LD1 F0_11_5 ( .D(\din[5][11] ), .G(n73), .Q(\q[5][11] ) );
    LD1 F0_4_13 ( .D(\din[13][4] ), .G(n73), .Q(\q[13][4] ) );
    LD1 F0_13_9 ( .D(\din[9][13] ), .G(n73), .Q(\q[9][13] ) );
    LD1 F0_3_1 ( .D(\din[1][3] ), .G(n73), .Q(\q[1][3] ) );
    LD1 F0_6_7 ( .D(\din[7][6] ), .G(n73), .Q(\q[7][6] ) );
    LD1 F0_11_12 ( .D(\din[12][11] ), .G(n73), .Q(\q[12][11] ) );
    LD1 F0_8_5 ( .D(\din[5][8] ), .G(n73), .Q(\q[5][8] ) );
    LD1 F0_5_12 ( .D(\din[12][5] ), .G(n73), .Q(\q[12][5] ) );
    LD1 F0_5_2 ( .D(\din[2][5] ), .G(n73), .Q(\q[2][5] ) );
    LD1 F0_2_1 ( .D(\din[1][2] ), .G(n73), .Q(\q[1][2] ) );
    LD1 F0_0_15 ( .D(\din[15][0] ), .G(n73), .Q(\q[15][0] ) );
    LD1 F0_14_12 ( .D(\din[12][14] ), .G(n73), .Q(\q[12][14] ) );
    LD1 F0_0_12 ( .D(\din[12][0] ), .G(n73), .Q(\q[12][0] ) );
    LD1 F0_12_0 ( .D(\din[0][12] ), .G(n73), .Q(\q[0][12] ) );
    LD1 F0_2_8 ( .D(\din[8][2] ), .G(n73), .Q(\q[8][2] ) );
    LD1 F0_0_4 ( .D(\din[4][0] ), .G(n73), .Q(\q[4][0] ) );
    LD1 F0_0_3 ( .D(\din[3][0] ), .G(n73), .Q(\q[3][0] ) );
    LD1 F0_13_0 ( .D(\din[0][13] ), .G(n73), .Q(\q[0][13] ) );
    LD1 F0_4_2 ( .D(\din[2][4] ), .G(n73), .Q(\q[2][4] ) );
    LD1 F0_3_8 ( .D(\din[8][3] ), .G(n73), .Q(\q[8][3] ) );
    LD1 F0_9_5 ( .D(\din[5][9] ), .G(n73), .Q(\q[5][9] ) );
    LD1 F0_1_13 ( .D(\din[13][1] ), .G(n73), .Q(\q[13][1] ) );
    LD1 F0_1_4 ( .D(\din[4][1] ), .G(n73), .Q(\q[4][1] ) );
    LD1 F0_15_13 ( .D(\din[13][15] ), .G(n73), .Q(\q[13][15] ) );
    LD1 F0_5_10 ( .D(\din[10][5] ), .G(n73), .Q(\q[10][5] ) );
    LD1 F0_11_10 ( .D(\din[10][11] ), .G(n73), .Q(\q[10][11] ) );
    LD1 F0_6_5 ( .D(\din[5][6] ), .G(n73), .Q(\q[5][6] ) );
    LD1 F0_3_15 ( .D(\din[15][3] ), .G(n73), .Q(\q[15][3] ) );
    LD1 F0_3_3 ( .D(\din[3][3] ), .G(n73), .Q(\q[3][3] ) );
    LD1 F0_11_7 ( .D(\din[7][11] ), .G(n73), .Q(\q[7][11] ) );
    LD1 F0_9_13 ( .D(\din[13][9] ), .G(n73), .Q(\q[13][9] ) );
    LD1 F0_14_1 ( .D(\din[1][14] ), .G(n73), .Q(\q[1][14] ) );
    LD1 F0_4_9 ( .D(\din[9][4] ), .G(n73), .Q(\q[9][4] ) );
    LD1 F0_4_11 ( .D(\din[11][4] ), .G(n73), .Q(\q[11][4] ) );
    LD1 F0_10_11 ( .D(\din[11][10] ), .G(n73), .Q(\q[11][10] ) );
    LD1 F0_7_5 ( .D(\din[5][7] ), .G(n73), .Q(\q[5][7] ) );
    LD1 F0_15_1 ( .D(\din[1][15] ), .G(n73), .Q(\q[1][15] ) );
    LD1 F0_10_7 ( .D(\din[7][10] ), .G(n73), .Q(\q[7][10] ) );
    LD1 F0_5_9 ( .D(\din[9][5] ), .G(n73), .Q(\q[9][5] ) );
    LD1 F0_2_3 ( .D(\din[3][2] ), .G(n73), .Q(\q[3][2] ) );
    LD1 F0_8_12 ( .D(\din[12][8] ), .G(n73), .Q(\q[12][8] ) );
    LD1 F0_2_14 ( .D(\din[14][2] ), .G(n73), .Q(\q[14][2] ) );
    LD1 F0_15_11 ( .D(\din[11][15] ), .G(n73), .Q(\q[11][15] ) );
    LD1 F0_13_2 ( .D(\din[2][13] ), .G(n73), .Q(\q[2][13] ) );
    LD1 F0_9_7 ( .D(\din[7][9] ), .G(n73), .Q(\q[7][9] ) );
    LD1 F0_14_8 ( .D(\din[8][14] ), .G(n73), .Q(\q[8][14] ) );
    LD1 F0_13_14 ( .D(\din[14][13] ), .G(n73), .Q(\q[14][13] ) );
    LD1 F0_4_0 ( .D(\din[0][4] ), .G(n73), .Q(\q[0][4] ) );
    LD1 F0_1_11 ( .D(\din[11][1] ), .G(n73), .Q(\q[11][1] ) );
    LD1 F0_0_2 ( .D(\din[2][0] ), .G(n73), .Q(\q[2][0] ) );
    LD1 F0_7_14 ( .D(\din[14][7] ), .G(n73), .Q(\q[14][7] ) );
    LD1 F0_12_2 ( .D(\din[2][12] ), .G(n73), .Q(\q[2][12] ) );
    LD1 F0_1_6 ( .D(\din[6][1] ), .G(n73), .Q(\q[6][1] ) );
    LD1 F0_14_10 ( .D(\din[10][14] ), .G(n73), .Q(\q[10][14] ) );
    LD1 F0_5_0 ( .D(\din[0][5] ), .G(n73), .Q(\q[0][5] ) );
    LD1 F0_15_8 ( .D(\din[8][15] ), .G(n73), .Q(\q[8][15] ) );
    LD1 F0_12_15 ( .D(\din[15][12] ), .G(n73), .Q(\q[15][12] ) );
    LD1 F0_8_7 ( .D(\din[7][8] ), .G(n73), .Q(\q[7][8] ) );
    LD1 F0_6_15 ( .D(\din[15][6] ), .G(n73), .Q(\q[15][6] ) );
    LD1 F0_12_12 ( .D(\din[12][12] ), .G(n73), .Q(\q[12][12] ) );
    LD1 F0_12_5 ( .D(\din[5][12] ), .G(n73), .Q(\q[5][12] ) );
    LD1 F0_8_0 ( .D(\din[0][8] ), .G(n73), .Q(\q[0][8] ) );
    LD1 F0_6_12 ( .D(\din[12][6] ), .G(n73), .Q(\q[12][6] ) );
    LD1 F0_10_9 ( .D(\din[9][10] ), .G(n73), .Q(\q[9][10] ) );
    LD1 F0_5_7 ( .D(\din[7][5] ), .G(n73), .Q(\q[7][5] ) );
    LD1 F0_0_10 ( .D(\din[10][0] ), .G(n73), .Q(\q[10][0] ) );
    LD1 F0_0_6 ( .D(\din[6][0] ), .G(n73), .Q(\q[6][0] ) );
    LD1 F0_13_5 ( .D(\din[5][13] ), .G(n73), .Q(\q[5][13] ) );
    LD1 F0_11_9 ( .D(\din[9][11] ), .G(n73), .Q(\q[9][11] ) );
    LD1 F0_7_13 ( .D(\din[13][7] ), .G(n73), .Q(\q[13][7] ) );
    LD1 F0_1_1 ( .D(\din[1][1] ), .G(n73), .Q(\q[1][1] ) );
    LD1 F0_13_13 ( .D(\din[13][13] ), .G(n73), .Q(\q[13][13] ) );
    LD1 F0_9_0 ( .D(\din[0][9] ), .G(n73), .Q(\q[0][9] ) );
    LD1 F0_4_7 ( .D(\din[7][4] ), .G(n73), .Q(\q[7][4] ) );
    LD1 F0_8_15 ( .D(\din[15][8] ), .G(n73), .Q(\q[15][8] ) );
    LD1 F0_8_9 ( .D(\din[9][8] ), .G(n73), .Q(\q[9][8] ) );
    LD1 F0_7_2 ( .D(\din[2][7] ), .G(n73), .Q(\q[2][7] ) );
    LD1 F0_2_13 ( .D(\din[13][2] ), .G(n73), .Q(\q[13][2] ) );
    LD1 F0_2_4 ( .D(\din[4][2] ), .G(n73), .Q(\q[4][2] ) );
    LD1 F0_10_0 ( .D(\din[0][10] ), .G(n73), .Q(\q[0][10] ) );
    LD1 F0_15_6 ( .D(\din[6][15] ), .G(n73), .Q(\q[6][15] ) );
    LD1 F0_3_4 ( .D(\din[4][3] ), .G(n73), .Q(\q[4][3] ) );
    LD1 F0_6_2 ( .D(\din[2][6] ), .G(n73), .Q(\q[2][6] ) );
    LD1 F0_14_6 ( .D(\din[6][14] ), .G(n73), .Q(\q[6][14] ) );
    LD1 F0_11_0 ( .D(\din[0][11] ), .G(n73), .Q(\q[0][11] ) );
    LD1 F0_9_14 ( .D(\din[14][9] ), .G(n73), .Q(\q[14][9] ) );
    LD1 F0_3_12 ( .D(\din[12][3] ), .G(n73), .Q(\q[12][3] ) );
    LD1 F0_9_9 ( .D(\din[9][9] ), .G(n73), .Q(\q[9][9] ) );
    LD1 F0_9_1 ( .D(\din[1][9] ), .G(n73), .Q(\q[1][9] ) );
    LD1 F0_13_4 ( .D(\din[4][13] ), .G(n73), .Q(\q[4][13] ) );
    LD1 F0_1_8 ( .D(\din[8][1] ), .G(n73), .Q(\q[8][1] ) );
    LD1 F0_1_0 ( .D(\din[0][1] ), .G(n73), .Q(\q[0][1] ) );
    LD1 F0_0_8 ( .D(\din[8][0] ), .G(n73), .Q(\q[8][0] ) );
    LD1 F0_11_8 ( .D(\din[8][11] ), .G(n73), .Q(\q[8][11] ) );
    LD1 F0_13_12 ( .D(\din[12][13] ), .G(n73), .Q(\q[12][13] ) );
    LD1 F0_7_12 ( .D(\din[12][7] ), .G(n73), .Q(\q[12][7] ) );
    LD1 F0_12_4 ( .D(\din[4][12] ), .G(n73), .Q(\q[4][12] ) );
    LD1 F0_4_6 ( .D(\din[6][4] ), .G(n73), .Q(\q[6][4] ) );
    LD1 F0_5_6 ( .D(\din[6][5] ), .G(n73), .Q(\q[6][5] ) );
    LD1 F0_10_8 ( .D(\din[8][10] ), .G(n73), .Q(\q[8][10] ) );
    LD1 F0_0_1 ( .D(\din[1][0] ), .G(n73), .Q(\q[1][0] ) );
    LD1 F0_12_13 ( .D(\din[13][12] ), .G(n73), .Q(\q[13][12] ) );
    LD1 F0_9_8 ( .D(\din[8][9] ), .G(n73), .Q(\q[8][9] ) );
    LD1 F0_8_1 ( .D(\din[1][8] ), .G(n73), .Q(\q[1][8] ) );
    LD1 F0_6_13 ( .D(\din[13][6] ), .G(n73), .Q(\q[13][6] ) );
    LD1 F0_6_3 ( .D(\din[3][6] ), .G(n73), .Q(\q[3][6] ) );
    LD1 F0_14_7 ( .D(\din[7][14] ), .G(n73), .Q(\q[7][14] ) );
    LD1 F0_11_1 ( .D(\din[1][11] ), .G(n73), .Q(\q[1][11] ) );
    LD1 F0_9_15 ( .D(\din[15][9] ), .G(n73), .Q(\q[15][9] ) );
    LD1 F0_3_13 ( .D(\din[13][3] ), .G(n73), .Q(\q[13][3] ) );
    LD1 F0_3_5 ( .D(\din[5][3] ), .G(n73), .Q(\q[5][3] ) );
    LD1 F0_7_3 ( .D(\din[3][7] ), .G(n73), .Q(\q[3][7] ) );
    LD1 F0_2_5 ( .D(\din[5][2] ), .G(n73), .Q(\q[5][2] ) );
    LD1 F0_1_9 ( .D(\din[9][1] ), .G(n73), .Q(\q[9][1] ) );
    LD1 F0_15_7 ( .D(\din[7][15] ), .G(n73), .Q(\q[7][15] ) );
    LD1 F0_10_1 ( .D(\din[1][10] ), .G(n73), .Q(\q[1][10] ) );
    LD1 F0_8_14 ( .D(\din[14][8] ), .G(n73), .Q(\q[14][8] ) );
    LD1 F0_8_8 ( .D(\din[8][8] ), .G(n73), .Q(\q[8][8] ) );
    LD1 F0_8_13 ( .D(\din[13][8] ), .G(n73), .Q(\q[13][8] ) );
    LD1 F0_4_10 ( .D(\din[10][4] ), .G(n73), .Q(\q[10][4] ) );
    LD1 F0_2_15 ( .D(\din[15][2] ), .G(n73), .Q(\q[15][2] ) );
    LD1 F0_2_12 ( .D(\din[12][2] ), .G(n73), .Q(\q[12][2] ) );
    LD1 F0_10_10 ( .D(\din[10][10] ), .G(n73), .Q(\q[10][10] ) );
    LD1 F0_15_0 ( .D(\din[0][15] ), .G(n73), .Q(\q[0][15] ) );
    LD1 F0_7_4 ( .D(\din[4][7] ), .G(n73), .Q(\q[4][7] ) );
    LD1 F0_5_8 ( .D(\din[8][5] ), .G(n73), .Q(\q[8][5] ) );
    LD1 F0_2_2 ( .D(\din[2][2] ), .G(n73), .Q(\q[2][2] ) );
    LD1 F0_10_6 ( .D(\din[6][10] ), .G(n73), .Q(\q[6][10] ) );
    LD1 F0_6_4 ( .D(\din[4][6] ), .G(n73), .Q(\q[4][6] ) );
    LD1 F0_3_14 ( .D(\din[14][3] ), .G(n73), .Q(\q[14][3] ) );
    LD1 F0_3_2 ( .D(\din[2][3] ), .G(n73), .Q(\q[2][3] ) );
    LD1 F0_0_9 ( .D(\din[9][0] ), .G(n73), .Q(\q[9][0] ) );
    LD1 F0_11_6 ( .D(\din[6][11] ), .G(n73), .Q(\q[6][11] ) );
    LD1 F0_14_0 ( .D(\din[0][14] ), .G(n73), .Q(\q[0][14] ) );
    LD1 F0_9_12 ( .D(\din[12][9] ), .G(n73), .Q(\q[12][9] ) );
    LD1 F0_5_11 ( .D(\din[11][5] ), .G(n73), .Q(\q[11][5] ) );
    LD1 F0_11_11 ( .D(\din[11][11] ), .G(n73), .Q(\q[11][11] ) );
    LD1 F0_12_14 ( .D(\din[14][12] ), .G(n73), .Q(\q[14][12] ) );
    LD1 F0_8_6 ( .D(\din[6][8] ), .G(n73), .Q(\q[6][8] ) );
    LD1 F0_14_11 ( .D(\din[11][14] ), .G(n73), .Q(\q[11][14] ) );
    LD1 F0_12_3 ( .D(\din[3][12] ), .G(n73), .Q(\q[3][12] ) );
    LD1 F0_6_14 ( .D(\din[14][6] ), .G(n73), .Q(\q[14][6] ) );
    LD1 F0_4_8 ( .D(\din[8][4] ), .G(n73), .Q(\q[8][4] ) );
    LD1 F0_15_9 ( .D(\din[9][15] ), .G(n73), .Q(\q[9][15] ) );
    LD1 F0_5_1 ( .D(\din[1][5] ), .G(n73), .Q(\q[1][5] ) );
    LD1 F0_14_9 ( .D(\din[9][14] ), .G(n73), .Q(\q[9][14] ) );
    LD1 F0_13_3 ( .D(\din[3][13] ), .G(n73), .Q(\q[3][13] ) );
    LD1 F0_13_15 ( .D(\din[15][13] ), .G(n73), .Q(\q[15][13] ) );
    LD1 F0_7_15 ( .D(\din[15][7] ), .G(n73), .Q(\q[15][7] ) );
    LD1 F0_4_1 ( .D(\din[1][4] ), .G(n73), .Q(\q[1][4] ) );
    LD1 F0_0_11 ( .D(\din[11][0] ), .G(n73), .Q(\q[11][0] ) );
    LD1 F0_0_7 ( .D(\din[7][0] ), .G(n73), .Q(\q[7][0] ) );
    LD1 F0_0_0 ( .D(\din[0][0] ), .G(n73), .Q(\q[0][0] ) );
    LD1 F0_1_7 ( .D(\din[7][1] ), .G(n73), .Q(\q[7][1] ) );
    LD1 F0_15_10 ( .D(\din[10][15] ), .G(n73), .Q(\q[10][15] ) );
    LD1 F0_9_6 ( .D(\din[6][9] ), .G(n73), .Q(\q[6][9] ) );
    LD1 F0_1_10 ( .D(\din[10][1] ), .G(n73), .Q(\q[10][1] ) );
    NR2 U72 ( .A(n91), .B(wr_n), .Z(\wren[6] ) );
    NR2 U73 ( .A(n92), .B(wr_n), .Z(\wren[1] ) );
    NR2 U74 ( .A(n93), .B(wr_n), .Z(\wren[8] ) );
    NR2 U75 ( .A(n95), .B(wr_n), .Z(\wren[10] ) );
    NR2 U76 ( .A(n96), .B(wr_n), .Z(\wren[0] ) );
    NR2 U77 ( .A(n97), .B(wr_n), .Z(\wren[11] ) );
    NR2 U78 ( .A(n98), .B(wr_n), .Z(\wren[9] ) );
    NR2 U79 ( .A(n99), .B(wr_n), .Z(\wren[7] ) );
    NR2 U80 ( .A(n100), .B(wr_n), .Z(\wren[14] ) );
    NR2 U81 ( .A(n101), .B(wr_n), .Z(\wren[5] ) );
    NR2 U82 ( .A(n102), .B(wr_n), .Z(\wren[2] ) );
    NR2 U83 ( .A(n103), .B(wr_n), .Z(\wren[13] ) );
    NR2 U84 ( .A(n104), .B(wr_n), .Z(\wren[3] ) );
    NR2 U85 ( .A(n105), .B(wr_n), .Z(\wren[12] ) );
    NR2 U86 ( .A(n106), .B(wr_n), .Z(\wren[15] ) );
    NR2 U87 ( .A(n107), .B(wr_n), .Z(\wren[4] ) );
    IV U88 ( .A(clk), .Z(n73) );
    IV U89 ( .A(wr_addr[9]), .Z(n98) );
    IV U90 ( .A(wr_addr[8]), .Z(n93) );
    IV U91 ( .A(wr_addr[7]), .Z(n99) );
    IV U92 ( .A(wr_addr[6]), .Z(n91) );
    IV U93 ( .A(wr_addr[5]), .Z(n101) );
    IV U94 ( .A(wr_addr[4]), .Z(n107) );
    IV U95 ( .A(wr_addr[3]), .Z(n104) );
    IV U96 ( .A(wr_addr[2]), .Z(n102) );
    IV U97 ( .A(wr_addr[1]), .Z(n92) );
    IV U98 ( .A(wr_addr[15]), .Z(n106) );
    IV U99 ( .A(wr_addr[14]), .Z(n100) );
    IV U100 ( .A(wr_addr[13]), .Z(n103) );
    IV U101 ( .A(wr_addr[12]), .Z(n105) );
    IV U102 ( .A(wr_addr[11]), .Z(n97) );
    IV U103 ( .A(wr_addr[10]), .Z(n95) );
    IV U104 ( .A(wr_addr[0]), .Z(n96) );
endmodule


module fifo_DW_ram_r_w_s_lat_32_16_0 ( clk, cs_n, wr_n, rd_addr, wr_addr, 
    data_in, data_out );
output [31:0] data_out;
input  [3:0] rd_addr;
input  [3:0] wr_addr;
input  [31:0] data_in;
input  clk, cs_n, wr_n;
    wire \addr_dec[13] , \addr_dec[15] , \addr_dec[11] , \addr_dec[4] , 
        \addr_dec[0] , \addr_dec[9] , \addr_dec[2] , \addr_dec[6] , 
        \addr_dec[7] , \addr_dec[3] , \addr_dec[1] , \addr_dec[8] , 
        \addr_dec[5] , \addr_dec[10] , \addr_dec[14] , \addr_dec[12] , n110, 
        n144, n145, n146, n147, n148, n149, n150, n151, n152, n153;
    fifo_DW_MEM_R_W_S_LAT_16_16_1 M0_2 ( .clk(clk), .wr_n(wr_n), .rd_addr(
        rd_addr), .wr_addr({\addr_dec[15] , \addr_dec[14] , \addr_dec[13] , 
        \addr_dec[12] , \addr_dec[11] , \addr_dec[10] , \addr_dec[9] , 
        \addr_dec[8] , \addr_dec[7] , \addr_dec[6] , \addr_dec[5] , 
        \addr_dec[4] , \addr_dec[3] , \addr_dec[2] , \addr_dec[1] , 
        \addr_dec[0] }), .data_in(data_in[15:0]), .data_out(data_out[15:0]) );
    fifo_DW_MEM_R_W_S_LAT_16_16_0 M0_1 ( .clk(clk), .wr_n(wr_n), .rd_addr(
        rd_addr), .wr_addr({\addr_dec[15] , \addr_dec[14] , \addr_dec[13] , 
        \addr_dec[12] , \addr_dec[11] , \addr_dec[10] , \addr_dec[9] , 
        \addr_dec[8] , \addr_dec[7] , \addr_dec[6] , \addr_dec[5] , 
        \addr_dec[4] , \addr_dec[3] , \addr_dec[2] , \addr_dec[1] , 
        \addr_dec[0] }), .data_in(data_in[31:16]), .data_out(data_out[31:16])
         );
    NR2 U60 ( .A(n110), .B(n144), .Z(\addr_dec[0] ) );
    NR2 U61 ( .A(n145), .B(n146), .Z(\addr_dec[10] ) );
    NR2 U62 ( .A(n147), .B(n146), .Z(\addr_dec[11] ) );
    NR2 U63 ( .A(n145), .B(n148), .Z(\addr_dec[12] ) );
    NR2 U64 ( .A(n147), .B(n148), .Z(\addr_dec[13] ) );
    NR2 U65 ( .A(n145), .B(n149), .Z(\addr_dec[14] ) );
    NR2 U66 ( .A(n147), .B(n149), .Z(\addr_dec[15] ) );
    NR2 U67 ( .A(n110), .B(n150), .Z(\addr_dec[1] ) );
    NR2 U68 ( .A(n144), .B(n146), .Z(\addr_dec[2] ) );
    NR2 U69 ( .A(n150), .B(n146), .Z(\addr_dec[3] ) );
    NR2 U70 ( .A(n144), .B(n148), .Z(\addr_dec[4] ) );
    NR2 U71 ( .A(n150), .B(n148), .Z(\addr_dec[5] ) );
    NR2 U72 ( .A(n149), .B(n144), .Z(\addr_dec[6] ) );
    NR2 U73 ( .A(n150), .B(n149), .Z(\addr_dec[7] ) );
    NR2 U74 ( .A(n110), .B(n145), .Z(\addr_dec[8] ) );
    NR2 U75 ( .A(n147), .B(n110), .Z(\addr_dec[9] ) );
    ND2 U76 ( .A(wr_addr[3]), .B(wr_addr[0]), .Z(n147) );
    ND2 U77 ( .A(n151), .B(n152), .Z(n110) );
    ND2 U78 ( .A(wr_addr[3]), .B(n153), .Z(n145) );
    IV U79 ( .A(wr_addr[2]), .Z(n151) );
    IV U80 ( .A(wr_addr[1]), .Z(n152) );
    OR2 U81 ( .A(n153), .B(wr_addr[3]), .Z(n150) );
    ND2 U82 ( .A(wr_addr[1]), .B(wr_addr[2]), .Z(n149) );
    ND3 U83 ( .A(n145), .B(n147), .C(n150), .Z(n144) );
    ND2 U84 ( .A(wr_addr[2]), .B(n152), .Z(n148) );
    ND2 U85 ( .A(wr_addr[1]), .B(n151), .Z(n146) );
    IV U86 ( .A(wr_addr[0]), .Z(n153) );
endmodule


module gray2bin_COUNT_WIDTH4_2 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U13 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U14 ( .A(gray_count[2]), .B(\gray_count[3] ), .Z(bin_count[2]) );
    EO U15 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module gray2bin_COUNT_WIDTH4_3 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U13 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U14 ( .A(gray_count[2]), .B(\gray_count[3] ), .Z(bin_count[2]) );
    EO U15 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module rs_flop_test_1 ( clk, reset_n, s, r, q_out, test_si, test_se );
input  [0:0] s;
output [0:0] q_out;
input  [0:0] r;
input  clk, reset_n, test_si, test_se;
    wire n112, n142, n143;
    FD1S \q_out_reg[0]  ( .D(n112), .CP(clk), .TI(test_si), .TE(test_se), .Q(
        q_out) );
    NR3 U14 ( .A(n142), .B(r), .C(n143), .Z(n112) );
    NR2 U15 ( .A(q_out), .B(s), .Z(n143) );
    IV U16 ( .A(reset_n), .Z(n142) );
endmodule


module gray_counter_WIDTH4_test_2 ( clk, reset, clear, enable, nxt_bin_count, 
    bin_count, gray_count, test_si, test_so, test_se );
output [3:0] nxt_bin_count;
output [3:0] gray_count;
output [3:0] bin_count;
input  clk, reset, clear, enable, test_si, test_se;
output test_so;
    wire n204, n208, n211, n215, n219, n223, n227, n231, n261, n262, n263, 
        n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
        n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
        n288, n289, n290, n291;
    assign gray_count[3] = test_so;
    FD1S \bin_count_reg[0]  ( .D(n211), .CP(clk), .TI(test_si), .TE(test_se), 
        .Q(bin_count[0]), .QN(n264) );
    FD1S \bin_count_reg[1]  ( .D(n215), .CP(clk), .TI(bin_count[0]), .TE(
        test_se), .Q(bin_count[1]), .QN(n263) );
    FD1S \bin_count_reg[2]  ( .D(n219), .CP(clk), .TI(bin_count[1]), .TE(
        test_se), .Q(bin_count[2]), .QN(n262) );
    FD1S \bin_count_reg[3]  ( .D(n223), .CP(clk), .TI(bin_count[2]), .TE(
        test_se), .Q(bin_count[3]), .QN(n261) );
    FD1S \prsnt_state_reg[0]  ( .D(n227), .CP(clk), .TI(bin_count[3]), .TE(
        test_se), .Q(gray_count[0]) );
    FD1S \prsnt_state_reg[3]  ( .D(n208), .CP(clk), .TI(gray_count[2]), .TE(
        test_se), .Q(test_so), .QN(n265) );
    FD1S \prsnt_state_reg[1]  ( .D(n231), .CP(clk), .TI(gray_count[0]), .TE(
        test_se), .Q(gray_count[1]), .QN(n266) );
    FD1S \prsnt_state_reg[2]  ( .D(n204), .CP(clk), .TI(gray_count[1]), .TE(
        test_se), .Q(gray_count[2]), .QN(n267) );
    AO7 U111 ( .A(n267), .B(n268), .C(n269), .Z(n204) );
    AO7 U112 ( .A(n265), .B(n268), .C(n270), .Z(n208) );
    EON1 U113 ( .A(n268), .B(n264), .C(n271), .D(nxt_bin_count[0]), .Z(n211)
         );
    AO7 U114 ( .A(n268), .B(n263), .C(n272), .Z(n215) );
    AO7 U115 ( .A(n268), .B(n262), .C(n273), .Z(n219) );
    AO7 U116 ( .A(n268), .B(n261), .C(n270), .Z(n223) );
    AO3 U117 ( .A(n274), .B(n272), .C(n275), .D(n276), .Z(n227) );
    AO7 U118 ( .A(n266), .B(n268), .C(n277), .Z(n231) );
    AO2 U119 ( .A(n265), .B(n267), .C(test_so), .D(gray_count[2]), .Z(n278) );
    AO2 U120 ( .A(n280), .B(n266), .C(n278), .D(gray_count[1]), .Z(n279) );
    EN U121 ( .A(gray_count[0]), .B(n279), .Z(n274) );
    EO1 U122 ( .A(test_so), .B(n282), .C(test_so), .D(n282), .Z(n281) );
    AO2 U123 ( .A(n280), .B(n284), .C(n278), .D(n285), .Z(n283) );
    IV U124 ( .A(enable), .Z(n286) );
    NR2 U125 ( .A(n286), .B(n274), .Z(n287) );
    ND2 U126 ( .A(n287), .B(n279), .Z(n285) );
    AO7 U127 ( .A(n287), .B(n279), .C(n285), .Z(n288) );
    AN2 U128 ( .A(reset), .B(enable), .Z(n271) );
    NR2 U129 ( .A(n283), .B(clear), .Z(nxt_bin_count[2]) );
    ND2 U130 ( .A(nxt_bin_count[2]), .B(n271), .Z(n273) );
    NR2 U131 ( .A(n288), .B(clear), .Z(nxt_bin_count[1]) );
    ND2 U132 ( .A(nxt_bin_count[1]), .B(n271), .Z(n272) );
    ND2 U133 ( .A(reset), .B(n286), .Z(n268) );
    AO1 U134 ( .A(n286), .B(n274), .C(clear), .D(n287), .Z(nxt_bin_count[0])
         );
    NR2 U135 ( .A(n281), .B(clear), .Z(nxt_bin_count[3]) );
    ND2 U136 ( .A(nxt_bin_count[3]), .B(n271), .Z(n270) );
    EO1 U137 ( .A(n289), .B(n288), .C(n272), .D(n290), .Z(n277) );
    EO1 U138 ( .A(n281), .B(n289), .C(n270), .D(n290), .Z(n269) );
    ND2 U139 ( .A(n284), .B(n278), .Z(n282) );
    IV U140 ( .A(n268), .Z(n291) );
    ND3 U141 ( .A(n288), .B(n271), .C(nxt_bin_count[0]), .Z(n275) );
    ND2 U142 ( .A(n291), .B(gray_count[0]), .Z(n276) );
    IV U143 ( .A(n283), .Z(n290) );
    IV U144 ( .A(n278), .Z(n280) );
    IV U145 ( .A(n285), .Z(n284) );
    IV U146 ( .A(n273), .Z(n289) );
endmodule


module push_ctrl_DEPTH16_counter_width4_almost_full_level8_test_1 ( push_clk, 
    reset_n, pop_count, push, push_full, almost_full, bin_count, push_count, 
    test_si, test_se );
input  [3:0] pop_count;
output [3:0] bin_count;
output [3:0] push_count;
input  push_clk, reset_n, push, test_si, test_se;
output push_full, almost_full;
    wire \pop_count_svd56[0] , \nxt_push_count[1] , \sync_pop_count[0] , 
        \sync_pop_count49[1] , count_enable, \sync_pop_count49[3] , 
        \sync_pop_count[2] , \nxt_push_count[3] , \pop_count_svd56[2] , 
        \sync_pop_countb[1] , \pop_count_svd[3] , counter_clear, 
        \pop_count_svdb[0] , \sync_pop_countb[3] , \pop_count_svd[1] , 
        \sync_pop_countb[2] , \pop_count_svd[0] , \pop_count_svd[2] , 
        \sync_pop_countb[0] , \sync_pop_count[3] , \nxt_push_count[2] , 
        make_full, internal_pop, \pop_count_svd56[3] , \sync_pop_count49[2] , 
        \sync_pop_count49[0] , \pop_count_svd56[1] , \nxt_push_count[0] , 
        \sync_pop_count[1] , n157, n158, n159, n160, n202, n292, n293, n294, 
        n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
        n307;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 ;
    gray2bin_COUNT_WIDTH4_3 synch1 ( .gray_count({\sync_pop_count[3] , 
        \sync_pop_count[2] , \sync_pop_count[1] , \sync_pop_count[0] }), 
        .bin_count({\sync_pop_countb[3] , \sync_pop_countb[2] , 
        \sync_pop_countb[1] , \sync_pop_countb[0] }) );
    gray2bin_COUNT_WIDTH4_2 synch2 ( .gray_count({\pop_count_svd[3] , 
        \pop_count_svd[2] , \pop_count_svd[1] , \pop_count_svd[0] }), 
        .bin_count({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, \pop_count_svdb[0] }) );
    rs_flop_test_1 full_flag ( .clk(push_clk), .reset_n(reset_n), .s(make_full
        ), .r(internal_pop), .q_out(push_full), .test_si(\sync_pop_count[3] ), 
        .test_se(test_se) );
    gray_counter_WIDTH4_test_2 push_counter ( .clk(push_clk), .reset(reset_n), 
        .clear(counter_clear), .enable(count_enable), .nxt_bin_count({
        \nxt_push_count[3] , \nxt_push_count[2] , \nxt_push_count[1] , 
        \nxt_push_count[0] }), .bin_count(bin_count), .gray_count(push_count), 
        .test_si(\pop_count_svd[3] ), .test_so(n202), .test_se(test_se) );
    FD1S \pop_count_svd_reg[0]  ( .D(\pop_count_svd56[0] ), .CP(push_clk), 
        .TI(test_si), .TE(test_se), .Q(\pop_count_svd[0] ) );
    FD1S \pop_count_svd_reg[1]  ( .D(\pop_count_svd56[1] ), .CP(push_clk), 
        .TI(\pop_count_svd[0] ), .TE(test_se), .Q(\pop_count_svd[1] ) );
    FD1S \pop_count_svd_reg[2]  ( .D(\pop_count_svd56[2] ), .CP(push_clk), 
        .TI(\pop_count_svd[1] ), .TE(test_se), .Q(\pop_count_svd[2] ) );
    FD1S \pop_count_svd_reg[3]  ( .D(\pop_count_svd56[3] ), .CP(push_clk), 
        .TI(\pop_count_svd[2] ), .TE(test_se), .Q(\pop_count_svd[3] ) );
    FD1S \sync_pop_count_reg[0]  ( .D(\sync_pop_count49[0] ), .CP(push_clk), 
        .TI(n202), .TE(test_se), .Q(\sync_pop_count[0] ), .QN(n160) );
    FD1S \sync_pop_count_reg[1]  ( .D(\sync_pop_count49[1] ), .CP(push_clk), 
        .TI(\sync_pop_count[0] ), .TE(test_se), .Q(\sync_pop_count[1] ), .QN(
        n159) );
    FD1S \sync_pop_count_reg[2]  ( .D(\sync_pop_count49[2] ), .CP(push_clk), 
        .TI(\sync_pop_count[1] ), .TE(test_se), .Q(\sync_pop_count[2] ), .QN(
        n158) );
    FD1S \sync_pop_count_reg[3]  ( .D(\sync_pop_count49[3] ), .CP(push_clk), 
        .TI(\sync_pop_count[2] ), .TE(test_se), .Q(\sync_pop_count[3] ), .QN(
        n157) );
    AN2 U71 ( .A(reset_n), .B(pop_count[3]), .Z(\sync_pop_count49[3] ) );
    AN2 U72 ( .A(pop_count[2]), .B(reset_n), .Z(\sync_pop_count49[2] ) );
    AN2 U73 ( .A(pop_count[1]), .B(reset_n), .Z(\sync_pop_count49[1] ) );
    AN2 U74 ( .A(pop_count[0]), .B(reset_n), .Z(\sync_pop_count49[0] ) );
    NR2 U75 ( .A(n292), .B(n157), .Z(\pop_count_svd56[3] ) );
    NR2 U76 ( .A(n292), .B(n158), .Z(\pop_count_svd56[2] ) );
    NR2 U77 ( .A(n292), .B(n159), .Z(\pop_count_svd56[1] ) );
    NR2 U78 ( .A(n292), .B(n160), .Z(\pop_count_svd56[0] ) );
    NR4 U79 ( .A(n293), .B(n294), .C(n295), .D(n296), .Z(make_full) );
    AN4 U80 ( .A(bin_count[2]), .B(bin_count[0]), .C(bin_count[1]), .D(
        bin_count[3]), .Z(counter_clear) );
    AN2 U81 ( .A(n297), .B(push), .Z(count_enable) );
    ND2 U82 ( .A(n298), .B(n297), .Z(almost_full) );
    EO1 U83 ( .A(bin_count[2]), .B(n300), .C(n301), .D(\sync_pop_countb[2] ), 
        .Z(n299) );
    IV U84 ( .A(reset_n), .Z(n292) );
    IV U85 ( .A(\sync_pop_countb[1] ), .Z(n302) );
    AO7 U86 ( .A(bin_count[1]), .B(n302), .C(n303), .Z(n301) );
    EO U87 ( .A(\sync_pop_countb[3] ), .B(\nxt_push_count[3] ), .Z(n293) );
    EO1 U88 ( .A(\sync_pop_countb[1] ), .B(\nxt_push_count[1] ), .C(
        \sync_pop_countb[1] ), .D(\nxt_push_count[1] ), .Z(n295) );
    EO1 U89 ( .A(\sync_pop_countb[2] ), .B(\nxt_push_count[2] ), .C(
        \sync_pop_countb[2] ), .D(\nxt_push_count[2] ), .Z(n296) );
    EO1 U90 ( .A(\sync_pop_countb[0] ), .B(\pop_count_svdb[0] ), .C(
        \sync_pop_countb[0] ), .D(\pop_count_svdb[0] ), .Z(internal_pop) );
    ND2 U91 ( .A(n304), .B(push), .Z(n294) );
    IV U92 ( .A(push_full), .Z(n297) );
    AO1 U93 ( .A(n302), .B(bin_count[1]), .C(bin_count[0]), .D(n306), .Z(n305)
         );
    ND2 U94 ( .A(\sync_pop_countb[2] ), .B(n301), .Z(n300) );
    EO1 U95 ( .A(\nxt_push_count[0] ), .B(n306), .C(\nxt_push_count[0] ), .D(
        n306), .Z(n304) );
    EO U96 ( .A(n299), .B(n307), .Z(n298) );
    EN U97 ( .A(bin_count[3]), .B(\sync_pop_countb[3] ), .Z(n307) );
    IV U98 ( .A(\sync_pop_countb[0] ), .Z(n306) );
    IV U99 ( .A(n305), .Z(n303) );
endmodule


module gray2bin_COUNT_WIDTH4_0 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U13 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U14 ( .A(gray_count[2]), .B(\gray_count[3] ), .Z(bin_count[2]) );
    EO U15 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module gray2bin_COUNT_WIDTH4_1 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U13 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U14 ( .A(gray_count[2]), .B(\gray_count[3] ), .Z(bin_count[2]) );
    EO U15 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module rs_flop_width1_reset_value1_test_1 ( clk, reset_n, s, r, q_out, test_si, 
    test_se );
input  [0:0] s;
output [0:0] q_out;
input  [0:0] r;
input  clk, reset_n, test_si, test_se;
    wire n91, n94;
    FD1S \q_out_reg[0]  ( .D(n91), .CP(clk), .TI(test_si), .TE(test_se), .Q(
        q_out) );
    AO7 U18 ( .A(r), .B(n94), .C(reset_n), .Z(n91) );
    NR2 U19 ( .A(q_out), .B(s), .Z(n94) );
endmodule


module gray_counter_WIDTH4_test_1 ( clk, reset, clear, enable, nxt_bin_count, 
    bin_count, gray_count, test_si, test_so, test_se );
output [3:0] nxt_bin_count;
output [3:0] gray_count;
output [3:0] bin_count;
input  clk, reset, clear, enable, test_si, test_se;
output test_so;
    wire n137, n141, n145, n149, n153, n157, n193, n197, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257;
    assign gray_count[3] = test_so;
    FD1S \bin_count_reg[0]  ( .D(n137), .CP(clk), .TI(test_si), .TE(test_se), 
        .Q(bin_count[0]), .QN(n230) );
    FD1S \bin_count_reg[1]  ( .D(n141), .CP(clk), .TI(bin_count[0]), .TE(
        test_se), .Q(bin_count[1]), .QN(n229) );
    FD1S \bin_count_reg[2]  ( .D(n145), .CP(clk), .TI(bin_count[1]), .TE(
        test_se), .Q(bin_count[2]), .QN(n228) );
    FD1S \bin_count_reg[3]  ( .D(n149), .CP(clk), .TI(bin_count[2]), .TE(
        test_se), .Q(bin_count[3]), .QN(n227) );
    FD1S \prsnt_state_reg[2]  ( .D(n193), .CP(clk), .TI(gray_count[1]), .TE(
        test_se), .Q(gray_count[2]) );
    FD1S \prsnt_state_reg[0]  ( .D(n153), .CP(clk), .TI(bin_count[3]), .TE(
        test_se), .Q(gray_count[0]) );
    FD1S \prsnt_state_reg[3]  ( .D(n197), .CP(clk), .TI(gray_count[2]), .TE(
        test_se), .Q(test_so), .QN(n231) );
    FD1S \prsnt_state_reg[1]  ( .D(n157), .CP(clk), .TI(gray_count[0]), .TE(
        test_se), .Q(gray_count[1]), .QN(n232) );
    EON1 U119 ( .A(n233), .B(n230), .C(n234), .D(nxt_bin_count[0]), .Z(n137)
         );
    AO7 U120 ( .A(n233), .B(n229), .C(n235), .Z(n141) );
    AO7 U121 ( .A(n233), .B(n228), .C(n236), .Z(n145) );
    AO7 U122 ( .A(n233), .B(n227), .C(n237), .Z(n149) );
    AO3 U123 ( .A(n238), .B(n235), .C(n239), .D(n240), .Z(n153) );
    AO7 U124 ( .A(n232), .B(n233), .C(n241), .Z(n157) );
    AO6 U125 ( .A(gray_count[2]), .B(n243), .C(n244), .Z(n242) );
    AO7 U126 ( .A(n231), .B(n233), .C(n237), .Z(n197) );
    EO1 U127 ( .A(test_so), .B(gray_count[2]), .C(test_so), .D(gray_count[2]), 
        .Z(n245) );
    AO2 U128 ( .A(n247), .B(n232), .C(n245), .D(gray_count[1]), .Z(n246) );
    EN U129 ( .A(gray_count[0]), .B(n246), .Z(n238) );
    EO1 U130 ( .A(test_so), .B(n249), .C(test_so), .D(n249), .Z(n248) );
    AO2 U131 ( .A(n247), .B(n251), .C(n245), .D(n252), .Z(n250) );
    IV U132 ( .A(enable), .Z(n253) );
    NR2 U133 ( .A(n253), .B(n238), .Z(n254) );
    ND2 U134 ( .A(n254), .B(n246), .Z(n252) );
    AO7 U135 ( .A(n254), .B(n246), .C(n252), .Z(n255) );
    ND2 U136 ( .A(reset), .B(n253), .Z(n233) );
    AN2 U137 ( .A(reset), .B(enable), .Z(n234) );
    NR2 U138 ( .A(n248), .B(clear), .Z(nxt_bin_count[3]) );
    NR2 U139 ( .A(n250), .B(clear), .Z(nxt_bin_count[2]) );
    ND2 U140 ( .A(nxt_bin_count[2]), .B(n234), .Z(n236) );
    ND2 U141 ( .A(nxt_bin_count[3]), .B(n234), .Z(n237) );
    NR2 U142 ( .A(n255), .B(clear), .Z(nxt_bin_count[1]) );
    ND2 U143 ( .A(nxt_bin_count[1]), .B(n234), .Z(n235) );
    AO1 U144 ( .A(n253), .B(n238), .C(clear), .D(n254), .Z(nxt_bin_count[0])
         );
    EON1 U145 ( .A(n237), .B(n256), .C(n257), .D(n248), .Z(n244) );
    EO1 U146 ( .A(n257), .B(n255), .C(n235), .D(n256), .Z(n241) );
    ND2 U147 ( .A(n251), .B(n245), .Z(n249) );
    IV U148 ( .A(n233), .Z(n243) );
    ND3 U149 ( .A(n255), .B(n234), .C(nxt_bin_count[0]), .Z(n239) );
    ND2 U150 ( .A(n243), .B(gray_count[0]), .Z(n240) );
    IV U151 ( .A(n250), .Z(n256) );
    IV U152 ( .A(n245), .Z(n247) );
    IV U153 ( .A(n252), .Z(n251) );
    IV U154 ( .A(n242), .Z(n193) );
    IV U155 ( .A(n236), .Z(n257) );
endmodule


module pop_ctrl_DEPTH16_counter_width4_almost_empty_level8_test_1 ( pop_clk, 
    reset_n, push_count, pop, pop_empty, almost_empty, bin_count, pop_count, 
    test_si, test_se );
input  [3:0] push_count;
output [3:0] bin_count;
output [3:0] pop_count;
input  pop_clk, reset_n, pop, test_si, test_se;
output pop_empty, almost_empty;
    wire \push_count_svd56[2] , \sync_push_count49[0] , \sync_push_count[0] , 
        count_enable, \sync_push_count[2] , \sync_push_count49[2] , 
        \push_count_svd56[0] , \nxt_pop_count[0] , \push_count_svd[0] , 
        \sync_push_countb[2] , counter_clear, \sync_push_countb[0] , 
        \push_count_svd[2] , \nxt_pop_count[2] , \push_count_svd[3] , 
        \nxt_pop_count[3] , \sync_push_countb[1] , \sync_push_countb[3] , 
        internal_push, \nxt_pop_count[1] , \push_count_svd[1] , 
        \sync_push_count49[3] , \push_count_svd56[1] , \sync_push_count[3] , 
        \sync_push_count[1] , \push_count_svdb[0] , make_empty, 
        \push_count_svd56[3] , \sync_push_count49[1] , n104, n105, n106, n107, 
        n109, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
        n137, n138, n139, n140, n141;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 ;
    gray2bin_COUNT_WIDTH4_1 synch1 ( .gray_count({\sync_push_count[3] , 
        \sync_push_count[2] , \sync_push_count[1] , \sync_push_count[0] }), 
        .bin_count({\sync_push_countb[3] , \sync_push_countb[2] , 
        \sync_push_countb[1] , \sync_push_countb[0] }) );
    gray2bin_COUNT_WIDTH4_0 synch2 ( .gray_count({\push_count_svd[3] , 
        \push_count_svd[2] , \push_count_svd[1] , \push_count_svd[0] }), 
        .bin_count({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, \push_count_svdb[0] }) );
    rs_flop_width1_reset_value1_test_1 empty_flag ( .clk(pop_clk), .reset_n(
        reset_n), .s(make_empty), .r(internal_push), .q_out(pop_empty), 
        .test_si(\sync_push_count[3] ), .test_se(test_se) );
    gray_counter_WIDTH4_test_1 push_counter ( .clk(pop_clk), .reset(reset_n), 
        .clear(counter_clear), .enable(count_enable), .nxt_bin_count({
        \nxt_pop_count[3] , \nxt_pop_count[2] , \nxt_pop_count[1] , 
        \nxt_pop_count[0] }), .bin_count(bin_count), .gray_count(pop_count), 
        .test_si(\push_count_svd[3] ), .test_so(n109), .test_se(test_se) );
    FD1S \push_count_svd_reg[0]  ( .D(\push_count_svd56[0] ), .CP(pop_clk), 
        .TI(test_si), .TE(test_se), .Q(\push_count_svd[0] ) );
    FD1S \push_count_svd_reg[1]  ( .D(\push_count_svd56[1] ), .CP(pop_clk), 
        .TI(\push_count_svd[0] ), .TE(test_se), .Q(\push_count_svd[1] ) );
    FD1S \push_count_svd_reg[2]  ( .D(\push_count_svd56[2] ), .CP(pop_clk), 
        .TI(\push_count_svd[1] ), .TE(test_se), .Q(\push_count_svd[2] ) );
    FD1S \push_count_svd_reg[3]  ( .D(\push_count_svd56[3] ), .CP(pop_clk), 
        .TI(\push_count_svd[2] ), .TE(test_se), .Q(\push_count_svd[3] ) );
    FD1S \sync_push_count_reg[0]  ( .D(\sync_push_count49[0] ), .CP(pop_clk), 
        .TI(n109), .TE(test_se), .Q(\sync_push_count[0] ), .QN(n107) );
    FD1S \sync_push_count_reg[1]  ( .D(\sync_push_count49[1] ), .CP(pop_clk), 
        .TI(\sync_push_count[0] ), .TE(test_se), .Q(\sync_push_count[1] ), 
        .QN(n106) );
    FD1S \sync_push_count_reg[2]  ( .D(\sync_push_count49[2] ), .CP(pop_clk), 
        .TI(\sync_push_count[1] ), .TE(test_se), .Q(\sync_push_count[2] ), 
        .QN(n105) );
    FD1S \sync_push_count_reg[3]  ( .D(\sync_push_count49[3] ), .CP(pop_clk), 
        .TI(\sync_push_count[2] ), .TE(test_se), .Q(\sync_push_count[3] ), 
        .QN(n104) );
    AN2 U71 ( .A(reset_n), .B(push_count[3]), .Z(\sync_push_count49[3] ) );
    AN2 U72 ( .A(push_count[2]), .B(reset_n), .Z(\sync_push_count49[2] ) );
    AN2 U73 ( .A(push_count[1]), .B(reset_n), .Z(\sync_push_count49[1] ) );
    AN2 U74 ( .A(push_count[0]), .B(reset_n), .Z(\sync_push_count49[0] ) );
    NR2 U75 ( .A(n126), .B(n104), .Z(\push_count_svd56[3] ) );
    NR2 U76 ( .A(n126), .B(n105), .Z(\push_count_svd56[2] ) );
    NR2 U77 ( .A(n126), .B(n106), .Z(\push_count_svd56[1] ) );
    NR2 U78 ( .A(n126), .B(n107), .Z(\push_count_svd56[0] ) );
    NR4 U79 ( .A(n127), .B(n128), .C(n129), .D(n130), .Z(make_empty) );
    AN4 U80 ( .A(bin_count[2]), .B(bin_count[0]), .C(bin_count[1]), .D(
        bin_count[3]), .Z(counter_clear) );
    AN2 U81 ( .A(n131), .B(pop), .Z(count_enable) );
    ND2 U82 ( .A(n132), .B(n131), .Z(almost_empty) );
    EO1 U83 ( .A(bin_count[2]), .B(n134), .C(n135), .D(\sync_push_countb[2] ), 
        .Z(n133) );
    IV U84 ( .A(reset_n), .Z(n126) );
    IV U85 ( .A(\sync_push_countb[1] ), .Z(n136) );
    AO7 U86 ( .A(bin_count[1]), .B(n136), .C(n137), .Z(n135) );
    EO U87 ( .A(\sync_push_countb[3] ), .B(\nxt_pop_count[3] ), .Z(n127) );
    EO1 U88 ( .A(\sync_push_countb[1] ), .B(\nxt_pop_count[1] ), .C(
        \sync_push_countb[1] ), .D(\nxt_pop_count[1] ), .Z(n129) );
    EO1 U89 ( .A(\sync_push_countb[2] ), .B(\nxt_pop_count[2] ), .C(
        \sync_push_countb[2] ), .D(\nxt_pop_count[2] ), .Z(n130) );
    EO1 U90 ( .A(\sync_push_countb[0] ), .B(\push_count_svdb[0] ), .C(
        \sync_push_countb[0] ), .D(\push_count_svdb[0] ), .Z(internal_push) );
    ND2 U91 ( .A(n138), .B(pop), .Z(n128) );
    IV U92 ( .A(pop_empty), .Z(n131) );
    AO1 U93 ( .A(n136), .B(bin_count[1]), .C(bin_count[0]), .D(n140), .Z(n139)
         );
    ND2 U94 ( .A(\sync_push_countb[2] ), .B(n135), .Z(n134) );
    EO1 U95 ( .A(\nxt_pop_count[0] ), .B(n140), .C(\nxt_pop_count[0] ), .D(
        n140), .Z(n138) );
    EO U96 ( .A(n133), .B(n141), .Z(n132) );
    EN U97 ( .A(bin_count[3]), .B(\sync_push_countb[3] ), .Z(n141) );
    IV U98 ( .A(\sync_push_countb[0] ), .Z(n140) );
    IV U99 ( .A(n139), .Z(n137) );
endmodule


module JTAG_BR ( CLOCKDR, SHIFTDR, TDI, TDO );
input  CLOCKDR, SHIFTDR, TDI;
output TDO;
    wire n8;
    FD1 U2 ( .D(n8), .CP(CLOCKDR), .Q(TDO) );
    AN2 U10 ( .A(SHIFTDR), .B(TDI), .Z(n8) );
endmodule


module JTAG_IR2 ( TDI, CLOCKIR, DI0, DI1, CLEAR0, CLEAR1, SET0, SET1, SHIFTIR, 
    UPDATEIR, TDO, DO0, DO1 );
input  TDI, CLOCKIR, DI0, DI1, CLEAR0, CLEAR1, SET0, SET1, SHIFTIR, UPDATEIR;
output TDO, DO0, DO1;
    wire n41, n42, n45, n53, n54, n55;
    FD3 OUT_BIT_1 ( .D(n45), .CP(UPDATEIR), .CD(CLEAR1), .SD(SET1), .Q(DO1) );
    FD1 SHADOW_BIT_1_1 ( .D(n42), .CP(CLOCKIR), .Q(n45) );
    FD3 OUT_BIT_0 ( .D(TDO), .CP(UPDATEIR), .CD(CLEAR0), .SD(SET0), .Q(DO0) );
    FD1 SHADOW_BIT_0_1 ( .D(n41), .CP(CLOCKIR), .Q(TDO) );
    AO2 U39 ( .A(DI1), .B(n54), .C(TDI), .D(SHIFTIR), .Z(n53) );
    AO2 U40 ( .A(DI0), .B(n54), .C(n45), .D(SHIFTIR), .Z(n55) );
    IV U41 ( .A(SHIFTIR), .Z(n54) );
    IV U42 ( .A(n53), .Z(n42) );
    IV U43 ( .A(n55), .Z(n41) );
endmodule


module JTAG_TAP ( TCK, TMS, TRST, CLOCKDR, CLOCKIR, ENABLE, RESET, SEL, 
    SHIFTDR, SHIFTIR, UPDATEDR, UPDATEIR );
input  TCK, TMS, TRST;
output CLOCKDR, CLOCKIR, ENABLE, RESET, SEL, SHIFTDR, SHIFTIR, UPDATEDR, 
    UPDATEIR;
    wire n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n111, 
        n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
        n124, n125;
    FD2 TAP_RESET_BAR ( .D(n96), .CP(n88), .CD(TRST), .Q(RESET) );
    FD2 TAP_SHIFTIR ( .D(n95), .CP(n88), .CD(TRST), .QN(SHIFTIR) );
    FD2 TAP_SHIFTDR ( .D(n94), .CP(n88), .CD(TRST), .QN(SHIFTDR) );
    FD2 TAP_ENABLE ( .D(n90), .CP(n88), .CD(TRST), .QN(ENABLE) );
    FD4 TAP_na ( .D(n91), .CP(TCK), .SD(TRST), .Q(n98), .QN(n111) );
    FD4 TAP_nd_SEL ( .D(n89), .CP(TCK), .SD(TRST), .Q(SEL), .QN(n112) );
    FD4 TAP_nc ( .D(n93), .CP(TCK), .SD(TRST), .Q(n97), .QN(n113) );
    FD4 TAP_nb ( .D(n92), .CP(TCK), .SD(TRST), .Q(n99), .QN(n114) );
    OR3 U105 ( .A(n115), .B(n113), .C(n114), .Z(n96) );
    AO4 U106 ( .A(n99), .B(n116), .C(n117), .D(n113), .Z(n93) );
    NR2 U107 ( .A(n115), .B(n118), .Z(UPDATEIR) );
    ND3 U108 ( .A(SEL), .B(n88), .C(n117), .Z(CLOCKIR) );
    IV U109 ( .A(TCK), .Z(n88) );
    ND2 U110 ( .A(n90), .B(n112), .Z(n94) );
    ND2 U111 ( .A(n90), .B(SEL), .Z(n95) );
    ND3 U112 ( .A(n88), .B(n112), .C(n117), .Z(CLOCKDR) );
    NR3 U113 ( .A(n111), .B(SEL), .C(n118), .Z(UPDATEDR) );
    AO3 U114 ( .A(n98), .B(SEL), .C(n97), .D(n120), .Z(n119) );
    AO1 U115 ( .A(n97), .B(SEL), .C(n114), .D(n111), .Z(n121) );
    AO6 U116 ( .A(n111), .B(n112), .C(n116), .Z(n122) );
    NR2 U117 ( .A(n99), .B(n113), .Z(n123) );
    ND2 U118 ( .A(SEL), .B(n98), .Z(n115) );
    NR2 U119 ( .A(n114), .B(n98), .Z(n117) );
    AN2 U120 ( .A(n117), .B(n113), .Z(n90) );
    ND3 U121 ( .A(n88), .B(n114), .C(n97), .Z(n118) );
    EO1 U122 ( .A(n124), .B(TMS), .C(n119), .D(TMS), .Z(n92) );
    AO2 U123 ( .A(n125), .B(n116), .C(n121), .D(TMS), .Z(n91) );
    EO1 U124 ( .A(n122), .B(n123), .C(SEL), .D(n123), .Z(n89) );
    ND2 U125 ( .A(n99), .B(n115), .Z(n120) );
    ND2 U126 ( .A(n97), .B(n120), .Z(n124) );
    ND2 U127 ( .A(n98), .B(n113), .Z(n125) );
    IV U128 ( .A(TMS), .Z(n116) );
endmodule


module JTAG_BSRINBOTH_0 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_1 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_2 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_3 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_4 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_5 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_6 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_7 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_8 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_9 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_10 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_11 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_12 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_13 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_14 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_15 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_16 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_17 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_18 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_19 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_20 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_21 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_22 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_23 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_24 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_25 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_26 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_27 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_28 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_29 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_30 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_31 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_32 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_33 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_34 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_35 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_36 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_37 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_38 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSRINBOTH_39 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n21, n22;
    FD1 SHADOW ( .D(n22), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n21) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n22) );
    EO1 U25 ( .A(n21), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_0 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_1 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_2 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_3 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_4 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_5 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_6 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_7 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_8 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_9 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_10 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_11 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_12 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_13 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_14 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_15 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_16 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_17 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_18 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_19 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_20 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_21 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_22 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_23 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_24 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_25 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_26 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_27 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_28 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_29 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_30 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_31 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_32 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_33 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_34 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module JTAG_BSROUTBOTH_35 ( TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11, TDO, 
    DO );
input  TDI, CLOCKDR, DI, SHIFTDR, UPDATEDR, MODE_11;
output TDO, DO;
    wire n23, n24;
    FD1 SHADOW ( .D(n24), .CP(CLOCKDR), .Q(TDO) );
    FD1 DATA_OUT ( .D(TDO), .CP(UPDATEDR), .QN(n23) );
    MUX21H U24 ( .A(DI), .B(TDI), .S(SHIFTDR), .Z(n24) );
    EO1 U25 ( .A(n23), .B(MODE_11), .C(DI), .D(MODE_11), .Z(DO) );
endmodule


module fifo ( push_clk, pop_clk, reset_n, push, pop, data_in, data_out, 
    pop_empty, push_full, almost_empty, almost_full, test_si1, test_si2, 
    test_se, jtag_tdo, jtag_tdi, jtag_tms, jtag_tck, jtag_trst );
input  [31:0] data_in;
output [31:0] data_out;
input  push_clk, pop_clk, reset_n, push, pop, test_si1, test_si2, test_se, 
    jtag_tdi, jtag_tms, jtag_tck, jtag_trst;
output pop_empty, push_full, almost_empty, almost_full, jtag_tdo;
    wire n493, n494, n496, n506, n510, n539, n550, n559, \dataout[6] , n519, 
        n543, n555, \push_count[2] , n502, n515, n535, \dataout[2] , n546, 
        n563, n504, n513, \rd_address[3] , \dataout[9] , \rd_address[1] , n537, 
        n557, \dataout[0] , n544, n497, n531, \push_count[0] , n532, n498, 
        n508, n517, n552, n541, n548, n561, n501, n521, n528, \dataout[4] , 
        \wr_address[0] , \dataout[25] , \dataout[16] , \pop_count[2] , n522, 
        n524, \dataout[21] , \dataout[12] , n565, \dataout[31] , \dataout[28] , 
        n562, \dataout[23] , \dataout[19] , \dataout[10] , n523, n526, 
        \pop_count[0] , n527, \pop_count[1] , \wr_address[2] , \dataout[27] , 
        \dataout[14] , n564, \wr_address[3] , \dataout[26] , \dataout[15] , 
        \dataout[22] , \dataout[18] , \dataout[11] , n525, \dataout[20] , 
        \dataout[13] , n529, \dataout[30] , \dataout[29] , \wr_address[1] , 
        \dataout[24] , \dataout[17] , \pop_count[3] , n495, n499, n500, n509, 
        n516, n520, n530, n533, \push_count[1] , n540, n553, n549, n505, n512, 
        n560, \dataout[5] , \rd_address[0] , \dataout[8] , n556, \dataout[1] , 
        n536, n545, n554, \dataout[3] , n534, n547, n503, n514, 
        \rd_address[2] , n511, n538, n57, n551, n558, \dataout[7] , n507, n518, 
        n542, \push_count[3] , n568, n567, n566, n313, n314, n315, n316, n317, 
        n318, n319, n320, n322, n324, n325, n326, n328, n330, n332, n334, n336, 
        n338, n340, n342, n344, n346, n348, n350, n352, n354, n356, n358, n360, 
        n362, n364, n366, n368, n370, n372, n374, n376, n378, n380, n382, n384, 
        n386, n388, n390, n392, n394, n396, n398, n400, n402, n404, n406, n408, 
        n410, n412, n414, n416, n418, n420, n422, n424, n426, n428, n430, n432, 
        n434, n436, n438, n440, n442, n444, n446, n448, n450, n452, n454, n456, 
        n458, n460, n462, n464, n466, n468, n470, n472, n474, n476, n477, n478, 
        n479, n481, n482, n483, n484, n485, n569, n570, n571, n572, n573, n574, 
        n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
        n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
        n599, n600, n601;
    tri jtag_tdo_wire;
    assign jtag_tdo = jtag_tdo_wire;
    fifo_DW_ram_r_w_s_lat_32_16_0 memory ( .clk(n493), .cs_n(1'b0), .wr_n(n57), 
        .rd_addr({\rd_address[3] , \rd_address[2] , \rd_address[1] , 
        \rd_address[0] }), .wr_addr({\wr_address[3] , \wr_address[2] , 
        \wr_address[1] , \wr_address[0] }), .data_in({n498, n499, n500, n501, 
        n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
        n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
        n526, n527, n528, n529}), .data_out({\dataout[31] , \dataout[30] , 
        \dataout[29] , \dataout[28] , \dataout[27] , \dataout[26] , 
        \dataout[25] , \dataout[24] , \dataout[23] , \dataout[22] , 
        \dataout[21] , \dataout[20] , \dataout[19] , \dataout[18] , 
        \dataout[17] , \dataout[16] , \dataout[15] , \dataout[14] , 
        \dataout[13] , \dataout[12] , \dataout[11] , \dataout[10] , 
        \dataout[9] , \dataout[8] , \dataout[7] , \dataout[6] , \dataout[5] , 
        \dataout[4] , \dataout[3] , \dataout[2] , \dataout[1] , \dataout[0] })
         );
    push_ctrl_DEPTH16_counter_width4_almost_full_level8_test_1 push_logic ( 
        .push_clk(n493), .reset_n(n495), .pop_count({\pop_count[3] , 
        \pop_count[2] , \pop_count[1] , \pop_count[0] }), .push(n496), 
        .push_full(n563), .almost_full(n565), .bin_count({\wr_address[3] , 
        \wr_address[2] , \wr_address[1] , \wr_address[0] }), .push_count({
        \push_count[3] , \push_count[2] , \push_count[1] , \push_count[0] }), 
        .test_si(n566), .test_se(n568) );
    pop_ctrl_DEPTH16_counter_width4_almost_empty_level8_test_1 pop_logic ( 
        .pop_clk(n494), .reset_n(n495), .push_count({\push_count[3] , 
        \push_count[2] , \push_count[1] , \push_count[0] }), .pop(n497), 
        .pop_empty(n562), .almost_empty(n564), .bin_count({\rd_address[3] , 
        \rd_address[2] , \rd_address[1] , \rd_address[0] }), .pop_count({
        \pop_count[3] , \pop_count[2] , \pop_count[1] , \pop_count[0] }), 
        .test_si(n567), .test_se(n568) );
    JTAG_BSRINBOTH_39 U154 ( .TDI(jtag_tdi), .CLOCKDR(n476), .DI(data_in[0]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n326), .DO(n529)
         );
    JTAG_BSRINBOTH_38 U155 ( .TDI(n326), .CLOCKDR(n476), .DI(data_in[1]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n328), .DO(n528)
         );
    JTAG_BSRINBOTH_37 U156 ( .TDI(n328), .CLOCKDR(n476), .DI(data_in[2]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n330), .DO(n527)
         );
    JTAG_BSRINBOTH_36 U157 ( .TDI(n330), .CLOCKDR(n476), .DI(data_in[3]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n332), .DO(n526)
         );
    JTAG_BSRINBOTH_35 U158 ( .TDI(n332), .CLOCKDR(n476), .DI(data_in[4]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n334), .DO(n525)
         );
    JTAG_BSRINBOTH_34 U159 ( .TDI(n334), .CLOCKDR(n476), .DI(data_in[5]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n336), .DO(n524)
         );
    JTAG_BSRINBOTH_33 U160 ( .TDI(n336), .CLOCKDR(n476), .DI(data_in[6]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n338), .DO(n523)
         );
    JTAG_BSRINBOTH_32 U161 ( .TDI(n338), .CLOCKDR(n476), .DI(data_in[7]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n340), .DO(n522)
         );
    JTAG_BSRINBOTH_31 U162 ( .TDI(n340), .CLOCKDR(n476), .DI(data_in[8]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n342), .DO(n521)
         );
    JTAG_BSRINBOTH_30 U163 ( .TDI(n342), .CLOCKDR(n476), .DI(data_in[9]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n344), .DO(n520)
         );
    JTAG_BSRINBOTH_29 U164 ( .TDI(n344), .CLOCKDR(n476), .DI(data_in[10]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n346), .DO(n519)
         );
    JTAG_BSRINBOTH_28 U165 ( .TDI(n346), .CLOCKDR(n476), .DI(data_in[11]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n348), .DO(n518)
         );
    JTAG_BSRINBOTH_27 U166 ( .TDI(n348), .CLOCKDR(n476), .DI(data_in[12]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n350), .DO(n517)
         );
    JTAG_BSRINBOTH_26 U167 ( .TDI(n350), .CLOCKDR(n476), .DI(data_in[13]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n352), .DO(n516)
         );
    JTAG_BSRINBOTH_25 U168 ( .TDI(n352), .CLOCKDR(n476), .DI(data_in[14]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n354), .DO(n515)
         );
    JTAG_BSRINBOTH_24 U169 ( .TDI(n354), .CLOCKDR(n476), .DI(data_in[15]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n356), .DO(n514)
         );
    JTAG_BSRINBOTH_23 U170 ( .TDI(n356), .CLOCKDR(n476), .DI(data_in[16]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n358), .DO(n513)
         );
    JTAG_BSRINBOTH_22 U171 ( .TDI(n358), .CLOCKDR(n476), .DI(data_in[17]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n360), .DO(n512)
         );
    JTAG_BSRINBOTH_21 U172 ( .TDI(n360), .CLOCKDR(n476), .DI(data_in[18]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n362), .DO(n511)
         );
    JTAG_BSRINBOTH_20 U173 ( .TDI(n362), .CLOCKDR(n476), .DI(data_in[19]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n364), .DO(n510)
         );
    JTAG_BSRINBOTH_19 U174 ( .TDI(n364), .CLOCKDR(n476), .DI(data_in[20]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n366), .DO(n509)
         );
    JTAG_BSRINBOTH_18 U175 ( .TDI(n366), .CLOCKDR(n476), .DI(data_in[21]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n368), .DO(n508)
         );
    JTAG_BSRINBOTH_17 U176 ( .TDI(n368), .CLOCKDR(n476), .DI(data_in[22]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n370), .DO(n507)
         );
    JTAG_BSRINBOTH_16 U177 ( .TDI(n370), .CLOCKDR(n476), .DI(data_in[23]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n372), .DO(n506)
         );
    JTAG_BSRINBOTH_15 U178 ( .TDI(n372), .CLOCKDR(n476), .DI(data_in[24]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n374), .DO(n505)
         );
    JTAG_BSRINBOTH_14 U179 ( .TDI(n374), .CLOCKDR(n476), .DI(data_in[25]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n376), .DO(n504)
         );
    JTAG_BSRINBOTH_13 U180 ( .TDI(n376), .CLOCKDR(n476), .DI(data_in[26]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n378), .DO(n503)
         );
    JTAG_BSRINBOTH_12 U181 ( .TDI(n378), .CLOCKDR(n476), .DI(data_in[27]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n380), .DO(n502)
         );
    JTAG_BSRINBOTH_11 U182 ( .TDI(n380), .CLOCKDR(n476), .DI(data_in[28]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n382), .DO(n501)
         );
    JTAG_BSRINBOTH_10 U183 ( .TDI(n382), .CLOCKDR(n476), .DI(data_in[29]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n384), .DO(n500)
         );
    JTAG_BSRINBOTH_9 U184 ( .TDI(n384), .CLOCKDR(n476), .DI(data_in[30]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n386), .DO(n499)
         );
    JTAG_BSRINBOTH_8 U185 ( .TDI(n386), .CLOCKDR(n476), .DI(data_in[31]), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n388), .DO(n498)
         );
    JTAG_BSRINBOTH_7 U186 ( .TDI(n388), .CLOCKDR(n476), .DI(pop), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n390), .DO(n497) );
    JTAG_BSRINBOTH_6 U187 ( .TDI(n390), .CLOCKDR(n476), .DI(pop_clk), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n392), .DO(n494)
         );
    JTAG_BSRINBOTH_5 U188 ( .TDI(n392), .CLOCKDR(n476), .DI(push), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n394), .DO(n496) );
    JTAG_BSRINBOTH_4 U189 ( .TDI(n394), .CLOCKDR(n476), .DI(push_clk), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n396), .DO(n493)
         );
    JTAG_BSRINBOTH_3 U190 ( .TDI(n396), .CLOCKDR(n476), .DI(reset_n), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n398), .DO(n495)
         );
    JTAG_BSRINBOTH_2 U191 ( .TDI(n398), .CLOCKDR(n476), .DI(test_se), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n400), .DO(n568)
         );
    JTAG_BSRINBOTH_1 U192 ( .TDI(n400), .CLOCKDR(n476), .DI(test_si1), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n402), .DO(n566)
         );
    JTAG_BSRINBOTH_0 BSR_IN_CELL ( .TDI(n402), .CLOCKDR(n476), .DI(test_si2), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n404), .DO(n567)
         );
    JTAG_BSROUTBOTH_35 U193 ( .TDI(n404), .CLOCKDR(n476), .DI(n564), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n406), .DO(almost_empty)
         );
    JTAG_BSROUTBOTH_34 U194 ( .TDI(n406), .CLOCKDR(n476), .DI(n565), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n408), .DO(almost_full)
         );
    JTAG_BSROUTBOTH_33 U195 ( .TDI(n408), .CLOCKDR(n476), .DI(n561), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n410), .DO(data_out[0])
         );
    JTAG_BSROUTBOTH_32 U196 ( .TDI(n410), .CLOCKDR(n476), .DI(n560), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n412), .DO(data_out[1])
         );
    JTAG_BSROUTBOTH_31 U197 ( .TDI(n412), .CLOCKDR(n476), .DI(n559), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n414), .DO(data_out[2])
         );
    JTAG_BSROUTBOTH_30 U198 ( .TDI(n414), .CLOCKDR(n476), .DI(n558), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n416), .DO(data_out[3])
         );
    JTAG_BSROUTBOTH_29 U199 ( .TDI(n416), .CLOCKDR(n476), .DI(n557), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n418), .DO(data_out[4])
         );
    JTAG_BSROUTBOTH_28 U200 ( .TDI(n418), .CLOCKDR(n476), .DI(n556), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n420), .DO(data_out[5])
         );
    JTAG_BSROUTBOTH_27 U201 ( .TDI(n420), .CLOCKDR(n476), .DI(n555), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n422), .DO(data_out[6])
         );
    JTAG_BSROUTBOTH_26 U202 ( .TDI(n422), .CLOCKDR(n476), .DI(n554), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n424), .DO(data_out[7])
         );
    JTAG_BSROUTBOTH_25 U203 ( .TDI(n424), .CLOCKDR(n476), .DI(n553), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n426), .DO(data_out[8])
         );
    JTAG_BSROUTBOTH_24 U204 ( .TDI(n426), .CLOCKDR(n476), .DI(n552), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n428), .DO(data_out[9])
         );
    JTAG_BSROUTBOTH_23 U205 ( .TDI(n428), .CLOCKDR(n476), .DI(n551), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n430), .DO(data_out[10])
         );
    JTAG_BSROUTBOTH_22 U206 ( .TDI(n430), .CLOCKDR(n476), .DI(n550), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n432), .DO(data_out[11])
         );
    JTAG_BSROUTBOTH_21 U207 ( .TDI(n432), .CLOCKDR(n476), .DI(n549), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n434), .DO(data_out[12])
         );
    JTAG_BSROUTBOTH_20 U208 ( .TDI(n434), .CLOCKDR(n476), .DI(n548), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n436), .DO(data_out[13])
         );
    JTAG_BSROUTBOTH_19 U209 ( .TDI(n436), .CLOCKDR(n476), .DI(n547), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n438), .DO(data_out[14])
         );
    JTAG_BSROUTBOTH_18 U210 ( .TDI(n438), .CLOCKDR(n476), .DI(n546), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n440), .DO(data_out[15])
         );
    JTAG_BSROUTBOTH_17 U211 ( .TDI(n440), .CLOCKDR(n476), .DI(n545), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n442), .DO(data_out[16])
         );
    JTAG_BSROUTBOTH_16 U212 ( .TDI(n442), .CLOCKDR(n476), .DI(n544), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n444), .DO(data_out[17])
         );
    JTAG_BSROUTBOTH_15 U213 ( .TDI(n444), .CLOCKDR(n476), .DI(n543), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n446), .DO(data_out[18])
         );
    JTAG_BSROUTBOTH_14 U214 ( .TDI(n446), .CLOCKDR(n476), .DI(n542), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n448), .DO(data_out[19])
         );
    JTAG_BSROUTBOTH_13 U215 ( .TDI(n448), .CLOCKDR(n476), .DI(n541), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n450), .DO(data_out[20])
         );
    JTAG_BSROUTBOTH_12 U216 ( .TDI(n450), .CLOCKDR(n476), .DI(n540), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n452), .DO(data_out[21])
         );
    JTAG_BSROUTBOTH_11 U217 ( .TDI(n452), .CLOCKDR(n476), .DI(n539), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n454), .DO(data_out[22])
         );
    JTAG_BSROUTBOTH_10 U218 ( .TDI(n454), .CLOCKDR(n476), .DI(n538), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n456), .DO(data_out[23])
         );
    JTAG_BSROUTBOTH_9 U219 ( .TDI(n456), .CLOCKDR(n476), .DI(n537), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n458), .DO(data_out[24])
         );
    JTAG_BSROUTBOTH_8 U220 ( .TDI(n458), .CLOCKDR(n476), .DI(n536), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n460), .DO(data_out[25])
         );
    JTAG_BSROUTBOTH_7 U221 ( .TDI(n460), .CLOCKDR(n476), .DI(n535), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n462), .DO(data_out[26])
         );
    JTAG_BSROUTBOTH_6 U222 ( .TDI(n462), .CLOCKDR(n476), .DI(n534), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n464), .DO(data_out[27])
         );
    JTAG_BSROUTBOTH_5 U223 ( .TDI(n464), .CLOCKDR(n476), .DI(n533), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n466), .DO(data_out[28])
         );
    JTAG_BSROUTBOTH_4 U224 ( .TDI(n466), .CLOCKDR(n476), .DI(n532), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n468), .DO(data_out[29])
         );
    JTAG_BSROUTBOTH_3 U225 ( .TDI(n468), .CLOCKDR(n476), .DI(n531), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n470), .DO(data_out[30])
         );
    JTAG_BSROUTBOTH_2 U226 ( .TDI(n470), .CLOCKDR(n476), .DI(n530), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n472), .DO(data_out[31])
         );
    JTAG_BSROUTBOTH_1 U227 ( .TDI(n472), .CLOCKDR(n476), .DI(n562), .SHIFTDR(
        n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n474), .DO(pop_empty) );
    JTAG_BSROUTBOTH_0 BSR_OUT_CELL ( .TDI(n474), .CLOCKDR(n476), .DI(n563), 
        .SHIFTDR(n477), .UPDATEDR(n324), .MODE_11(n325), .TDO(n317), .DO(
        push_full) );
    JTAG_BR JTAG_BYPASS_REG ( .CLOCKDR(n476), .SHIFTDR(n477), .TDI(jtag_tdi), 
        .TDO(n316) );
    JTAG_IR2 JTAG_IR ( .TDI(jtag_tdi), .CLOCKIR(n481), .DI0(1'b1), .DI1(1'b0), 
        .CLEAR0(1'b1), .CLEAR1(1'b1), .SET0(n485), .SET1(n485), .SHIFTIR(n482), 
        .UPDATEIR(n483), .TDO(n318), .DO0(n478), .DO1(n479) );
    JTAG_TAP JTAG_TAP_CONTROLLER ( .TCK(jtag_tck), .TMS(jtag_tms), .TRST(
        jtag_trst), .CLOCKDR(n476), .CLOCKIR(n481), .ENABLE(n322), .RESET(n484
        ), .SEL(n319), .SHIFTDR(n477), .SHIFTIR(n482), .UPDATEDR(n324), 
        .UPDATEIR(n483) );
    BTS4 U152 ( .A(n313), .E(n314), .Z(jtag_tdo_wire) );
    FD1 U153 ( .D(n320), .CP(n315), .Q(n313) );
    IV U232 ( .A(n496), .Z(n57) );
    NR2 U233 ( .A(n569), .B(n562), .Z(n530) );
    NR2 U234 ( .A(n570), .B(n562), .Z(n531) );
    NR2 U235 ( .A(n571), .B(n562), .Z(n532) );
    NR2 U236 ( .A(n572), .B(n562), .Z(n533) );
    NR2 U237 ( .A(n573), .B(n562), .Z(n534) );
    NR2 U238 ( .A(n574), .B(n562), .Z(n535) );
    NR2 U239 ( .A(n575), .B(n562), .Z(n536) );
    NR2 U240 ( .A(n576), .B(n562), .Z(n537) );
    NR2 U241 ( .A(n577), .B(n562), .Z(n538) );
    NR2 U242 ( .A(n578), .B(n562), .Z(n539) );
    NR2 U243 ( .A(n579), .B(n562), .Z(n540) );
    NR2 U244 ( .A(n580), .B(n562), .Z(n541) );
    NR2 U245 ( .A(n581), .B(n562), .Z(n542) );
    NR2 U246 ( .A(n582), .B(n562), .Z(n543) );
    NR2 U247 ( .A(n583), .B(n562), .Z(n544) );
    NR2 U248 ( .A(n584), .B(n562), .Z(n545) );
    NR2 U249 ( .A(n585), .B(n562), .Z(n546) );
    NR2 U250 ( .A(n586), .B(n562), .Z(n547) );
    NR2 U251 ( .A(n587), .B(n562), .Z(n548) );
    NR2 U252 ( .A(n588), .B(n562), .Z(n549) );
    NR2 U253 ( .A(n589), .B(n562), .Z(n550) );
    NR2 U254 ( .A(n590), .B(n562), .Z(n551) );
    NR2 U255 ( .A(n591), .B(n562), .Z(n552) );
    NR2 U256 ( .A(n592), .B(n562), .Z(n553) );
    NR2 U257 ( .A(n593), .B(n562), .Z(n554) );
    NR2 U258 ( .A(n594), .B(n562), .Z(n555) );
    NR2 U259 ( .A(n595), .B(n562), .Z(n556) );
    NR2 U260 ( .A(n596), .B(n562), .Z(n557) );
    NR2 U261 ( .A(n597), .B(n562), .Z(n558) );
    NR2 U262 ( .A(n598), .B(n562), .Z(n559) );
    NR2 U263 ( .A(n599), .B(n562), .Z(n560) );
    NR2 U264 ( .A(n600), .B(n562), .Z(n561) );
    AN2 U265 ( .A(jtag_trst), .B(n484), .Z(n485) );
    NR2 U266 ( .A(n478), .B(n479), .Z(n325) );
    IV U267 ( .A(jtag_tck), .Z(n315) );
    IV U268 ( .A(n322), .Z(n314) );
    MUX31L U269 ( .D0(n317), .D1(n316), .D2(n318), .A(n479), .B(n319), .Z(n601
        ) );
    IV U270 ( .A(n601), .Z(n320) );
    IV U271 ( .A(\dataout[0] ), .Z(n600) );
    IV U272 ( .A(\dataout[1] ), .Z(n599) );
    IV U273 ( .A(\dataout[2] ), .Z(n598) );
    IV U274 ( .A(\dataout[3] ), .Z(n597) );
    IV U275 ( .A(\dataout[4] ), .Z(n596) );
    IV U276 ( .A(\dataout[5] ), .Z(n595) );
    IV U277 ( .A(\dataout[6] ), .Z(n594) );
    IV U278 ( .A(\dataout[7] ), .Z(n593) );
    IV U279 ( .A(\dataout[8] ), .Z(n592) );
    IV U280 ( .A(\dataout[9] ), .Z(n591) );
    IV U281 ( .A(\dataout[10] ), .Z(n590) );
    IV U282 ( .A(\dataout[11] ), .Z(n589) );
    IV U283 ( .A(\dataout[12] ), .Z(n588) );
    IV U284 ( .A(\dataout[13] ), .Z(n587) );
    IV U285 ( .A(\dataout[14] ), .Z(n586) );
    IV U286 ( .A(\dataout[15] ), .Z(n585) );
    IV U287 ( .A(\dataout[16] ), .Z(n584) );
    IV U288 ( .A(\dataout[17] ), .Z(n583) );
    IV U289 ( .A(\dataout[18] ), .Z(n582) );
    IV U290 ( .A(\dataout[19] ), .Z(n581) );
    IV U291 ( .A(\dataout[20] ), .Z(n580) );
    IV U292 ( .A(\dataout[21] ), .Z(n579) );
    IV U293 ( .A(\dataout[22] ), .Z(n578) );
    IV U294 ( .A(\dataout[23] ), .Z(n577) );
    IV U295 ( .A(\dataout[24] ), .Z(n576) );
    IV U296 ( .A(\dataout[25] ), .Z(n575) );
    IV U297 ( .A(\dataout[26] ), .Z(n574) );
    IV U298 ( .A(\dataout[27] ), .Z(n573) );
    IV U299 ( .A(\dataout[28] ), .Z(n572) );
    IV U300 ( .A(\dataout[29] ), .Z(n571) );
    IV U301 ( .A(\dataout[30] ), .Z(n570) );
    IV U302 ( .A(\dataout[31] ), .Z(n569) );
endmodule

